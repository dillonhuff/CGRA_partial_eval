//Module: highImpedanceBit defined externally
//Module: pullresistor defined externally


module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule //corebit_and

module coreir_orr #(parameter width=1) (
  input [width-1:0] in,
  output out
);
  assign out = |in;

endmodule //coreir_orr

module corebit_mux (
  input in0,
  input in1,
  input sel,
  output out
);
  assign out = sel ? in1 : in0;

endmodule //corebit_mux

module coreir_xor #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 ^ in1;

endmodule //coreir_xor

module coreir_zext #(parameter width_in=1, parameter width_out=1) (
  input [width_in-1:0] in,
  output [width_out-1:0] out
);
  assign out = {{(width_out-width_in){1'b0}},in};

endmodule //coreir_zext

module coreir_or #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 | in1;

endmodule //coreir_or

module coreir_andr #(parameter width=1) (
  input [width-1:0] in,
  output out
);
  assign out = &in;

endmodule //coreir_andr

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule //coreir_eq

module corebit_concat (
  input in0,
  input in1,
  output [1:0] out
);
  assign out = {in0, in1};

endmodule //corebit_concat

module test_lut (
  input [7:0] cfg_a,
  input  cfg_clk,
  input [31:0] cfg_d,
  input  cfg_en,
  input  cfg_rst_n,
  input [15:0] op_a_in,
  input [15:0] op_b_in,
  input  op_c_in,
  output [15:0] res
);
  //All the connections
  assign res[0] = op_a_in[0];
  assign res[1] = op_a_in[1];
  assign res[10] = op_a_in[10];
  assign res[11] = op_a_in[11];
  assign res[12] = op_a_in[12];
  assign res[13] = op_a_in[13];
  assign res[14] = op_a_in[14];
  assign res[15] = op_a_in[15];
  assign res[2] = op_a_in[2];
  assign res[3] = op_a_in[3];
  assign res[4] = op_a_in[4];
  assign res[5] = op_a_in[5];
  assign res[6] = op_a_in[6];
  assign res[7] = op_a_in[7];
  assign res[8] = op_a_in[8];
  assign res[9] = op_a_in[9];

endmodule //test_lut

module corebit_tribuf (
  input in,
  input en,
  inout out
);
  assign out = en ? in : 1'bz;

endmodule //corebit_tribuf

module coreir_mux #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  input sel,
  output [width-1:0] out
);
  assign out = sel ? in1 : in0;

endmodule //coreir_mux

module coreir_add #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 + in1;

endmodule //coreir_add

module coreir_and #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 & in1;

endmodule //coreir_and

module corebit_or (
  input in0,
  input in1,
  output out
);
  assign out = in0 | in1;

endmodule //corebit_or

module reduce_or_U40 (
  input [7:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [7:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(8)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[7:0] = A[7:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U40

module corebit_wire (
  input in,
  output out
);
  assign out = in;

endmodule //corebit_wire

module coreir_not #(parameter width=1) (
  input [width-1:0] in,
  output [width-1:0] out
);
  assign out = ~in;

endmodule //coreir_not

module corebit_not (
  input in,
  output out
);
  assign out = ~in;

endmodule //corebit_not

module coreir_lshr #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 >> in1;

endmodule //coreir_lshr

module coreir_mul #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 * in1;

endmodule //coreir_mul

module corebit_term (
  input in
);


endmodule //corebit_term

module coreir_ashr #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = $signed(in0) >>> in1;

endmodule //coreir_ashr

module reduce_or_U30 (
  input [3:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [3:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(4)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[3:0] = A[3:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U30

module reduce_or_U37 (
  input [15:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [15:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(16)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[15:0] = A[15:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U37

module reduce_or_U29 (
  input [4:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [4:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(5)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[4:0] = A[4:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U29

module coreir_reg_arst #(parameter arst_posedge=1, parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input arst,
  input [width-1:0] in,
  output [width-1:0] out
);
reg [width-1:0] outReg;
wire real_rst;
assign real_rst = arst_posedge ? arst : ~arst;
wire real_clk;
assign real_clk = clk_posedge ? clk : ~clk;
always @(posedge real_clk, posedge real_rst) begin
  if (real_rst) outReg <= init;
  else outReg <= in;
end
assign out = outReg;

endmodule //coreir_reg_arst

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule //corebit_const

module __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__1 (
  input  cfg_clk,
  input  cfg_d,
  input  cfg_en,
  input  cfg_rst_n,
  input  data_in,
  output  debug_irq
);
  //Wire declarations for instance 'self__DOT__debug_irq__DOLLAR__bit_const_0' (Module corebit_const)
  wire  self__DOT__debug_irq__DOLLAR__bit_const_0__out;
  corebit_const #(.value(0)) self__DOT__debug_irq__DOLLAR__bit_const_0(
    .out(self__DOT__debug_irq__DOLLAR__bit_const_0__out)
  );

  //All the connections
  assign debug_irq = self__DOT__debug_irq__DOLLAR__bit_const_0__out;

endmodule //__DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__1

module add_U1 (
  input [15:0] A,
  input [15:0] B,
  output [16:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [16:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(17)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [15:0] extendB__in;
  wire [16:0] extendB__out;
  coreir_zext #(.width_in(16),.width_out(17)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_add)
  wire [16:0] op0__in0;
  wire [16:0] op0__in1;
  wire [16:0] op0__out;
  coreir_add #(.width(17)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[16:0] = extendA__out[16:0];
  assign extendB__in[15:0] = B[15:0];
  assign op0__in1[16:0] = extendB__out[16:0];
  assign Y[16:0] = op0__out[16:0];

endmodule //add_U1

module coreir_const #(parameter value=1, parameter width=1) (
  output [width-1:0] out
);
  assign out = value;

endmodule //coreir_const

module coreir_slice #(parameter hi=1, parameter lo=1, parameter width=1) (
  input [width-1:0] in,
  output [hi-lo-1:0] out
);
  assign out = in[hi-1:lo];

endmodule //coreir_slice

module coreir_ult #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 < in1;

endmodule //coreir_ult

module coreir_wrap (
  input in,
  output out
);
  assign out = in;

endmodule //coreir_wrap

module add_U11 (
  input [3:0] A,
  input [31:0] B,
  output [31:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [3:0] extendA__in;
  wire [31:0] extendA__out;
  coreir_zext #(.width_in(4),.width_out(32)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [31:0] extendB__in;
  wire [31:0] extendB__out;
  coreir_zext #(.width_in(32),.width_out(32)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_add)
  wire [31:0] op0__in0;
  wire [31:0] op0__in1;
  wire [31:0] op0__out;
  coreir_add #(.width(32)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[3:0] = A[3:0];
  assign op0__in0[31:0] = extendA__out[31:0];
  assign extendB__in[31:0] = B[31:0];
  assign op0__in1[31:0] = extendB__out[31:0];
  assign Y[31:0] = op0__out[31:0];

endmodule //add_U11

module eq_U18 (
  input [2:0] A,
  input [2:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [2:0] extendA__in;
  wire [2:0] extendA__out;
  coreir_zext #(.width_in(3),.width_out(3)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [2:0] extendB__in;
  wire [2:0] extendB__out;
  coreir_zext #(.width_in(3),.width_out(3)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [2:0] op0__in0;
  wire [2:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(3)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[2:0] = A[2:0];
  assign op0__in0[2:0] = extendA__out[2:0];
  assign extendB__in[2:0] = B[2:0];
  assign op0__in1[2:0] = extendB__out[2:0];
  assign Y[0] = op0__out;

endmodule //eq_U18

module corebit_ibuf (
  inout in,
  output out
);
  assign out = in;

endmodule //corebit_ibuf

module xor_U41 (
  input [15:0] A,
  input [15:0] B,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [15:0] extendB__in;
  wire [15:0] extendB__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_xor)
  wire [15:0] op0__in0;
  wire [15:0] op0__in1;
  wire [15:0] op0__out;
  coreir_xor #(.width(16)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[15:0] = extendA__out[15:0];
  assign extendB__in[15:0] = B[15:0];
  assign op0__in1[15:0] = extendB__out[15:0];
  assign Y[15:0] = op0__out[15:0];

endmodule //xor_U41

module not_U35 (
  input [15:0] A,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_not)
  wire [15:0] op0__in;
  wire [15:0] op0__out;
  coreir_not #(.width(16)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in[15:0] = extendA__out[15:0];
  assign Y[15:0] = op0__out[15:0];

endmodule //not_U35

module or_U6 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_or)
  wire [0:0] op0__in0;
  wire [0:0] op0__in1;
  wire [0:0] op0__out;
  coreir_or #(.width(1)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in0[0:0] = extendA__out[0:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[0:0] = extendB__out[0:0];
  assign Y[0:0] = op0__out[0:0];

endmodule //or_U6

module not_U14 (
  input [0:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_not)
  wire [0:0] op0__in;
  wire [0:0] op0__out;
  coreir_not #(.width(1)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in[0:0] = extendA__out[0:0];
  assign Y[0:0] = op0__out[0:0];

endmodule //not_U14

module test_debug_reg (
  input  cfg_clk,
  input [15:0] cfg_d,
  input  cfg_en,
  input  cfg_rst_n,
  input [15:0] data_in,
  output  debug_irq
);
  //Wire declarations for instance 'self__DOT__debug_irq__DOLLAR__bit_const_0' (Module corebit_const)
  wire  self__DOT__debug_irq__DOLLAR__bit_const_0__out;
  corebit_const #(.value(0)) self__DOT__debug_irq__DOLLAR__bit_const_0(
    .out(self__DOT__debug_irq__DOLLAR__bit_const_0__out)
  );

  //All the connections
  assign debug_irq = self__DOT__debug_irq__DOLLAR__bit_const_0__out;

endmodule //test_debug_reg

module corebit_xor (
  input in0,
  input in1,
  output out
);
  assign out = in0 ^ in1;

endmodule //corebit_xor

module eq_U17 (
  input [7:0] A,
  input [7:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [7:0] extendA__in;
  wire [7:0] extendA__out;
  coreir_zext #(.width_in(8),.width_out(8)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [7:0] extendB__in;
  wire [7:0] extendB__out;
  coreir_zext #(.width_in(8),.width_out(8)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [7:0] op0__in0;
  wire [7:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(8)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[7:0] = A[7:0];
  assign op0__in0[7:0] = extendA__out[7:0];
  assign extendB__in[7:0] = B[7:0];
  assign op0__in1[7:0] = extendB__out[7:0];
  assign Y[0] = op0__out;

endmodule //eq_U17

module eq_U32 (
  input [5:0] A,
  input [5:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [5:0] extendA__in;
  wire [5:0] extendA__out;
  coreir_zext #(.width_in(6),.width_out(6)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [5:0] extendB__in;
  wire [5:0] extendB__out;
  coreir_zext #(.width_in(6),.width_out(6)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [5:0] op0__in0;
  wire [5:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(6)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[5:0] = A[5:0];
  assign op0__in0[5:0] = extendA__out[5:0];
  assign extendB__in[5:0] = B[5:0];
  assign op0__in1[5:0] = extendB__out[5:0];
  assign Y[0] = op0__out;

endmodule //eq_U32

module lt_U20 (
  input [2:0] A,
  input [31:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [2:0] extendA__in;
  wire [31:0] extendA__out;
  coreir_zext #(.width_in(3),.width_out(32)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [31:0] extendB__in;
  wire [31:0] extendB__out;
  coreir_zext #(.width_in(32),.width_out(32)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_ult)
  wire [31:0] op0__in0;
  wire [31:0] op0__in1;
  wire  op0__out;
  coreir_ult #(.width(32)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[2:0] = A[2:0];
  assign op0__in0[31:0] = extendA__out[31:0];
  assign extendB__in[31:0] = B[31:0];
  assign op0__in1[31:0] = extendB__out[31:0];
  assign Y[0] = op0__out;

endmodule //lt_U20

module mul_U4 (
  input [16:0] A,
  input [16:0] B,
  output [33:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [16:0] extendA__in;
  wire [33:0] extendA__out;
  coreir_zext #(.width_in(17),.width_out(34)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [16:0] extendB__in;
  wire [33:0] extendB__out;
  coreir_zext #(.width_in(17),.width_out(34)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_mul)
  wire [33:0] op0__in0;
  wire [33:0] op0__in1;
  wire [33:0] op0__out;
  coreir_mul #(.width(34)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[16:0] = A[16:0];
  assign op0__in0[33:0] = extendA__out[33:0];
  assign extendB__in[16:0] = B[16:0];
  assign op0__in1[33:0] = extendB__out[33:0];
  assign Y[33:0] = op0__out[33:0];

endmodule //mul_U4

module sshr_U22 (
  input [15:0] A,
  input [3:0] B,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [3:0] extendB__in;
  wire [15:0] extendB__out;
  coreir_zext #(.width_in(4),.width_out(16)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_ashr)
  wire [15:0] op0__in0;
  wire [15:0] op0__in1;
  wire [15:0] op0__out;
  coreir_ashr #(.width(16)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //Wire declarations for instance 'slice0' (Module coreir_slice)
  wire [15:0] slice0__in;
  wire [15:0] slice0__out;
  coreir_slice #(.hi(16),.lo(0),.width(16)) slice0(
    .in(slice0__in),
    .out(slice0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[15:0] = extendA__out[15:0];
  assign extendB__in[3:0] = B[3:0];
  assign op0__in1[15:0] = extendB__out[15:0];
  assign slice0__in[15:0] = op0__out[15:0];
  assign Y[15:0] = slice0__out[15:0];

endmodule //sshr_U22

module shr_U21 (
  input [15:0] A,
  input [3:0] B,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [3:0] extendB__in;
  wire [15:0] extendB__out;
  coreir_zext #(.width_in(4),.width_out(16)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_lshr)
  wire [15:0] op0__in0;
  wire [15:0] op0__in1;
  wire [15:0] op0__out;
  coreir_lshr #(.width(16)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //Wire declarations for instance 'slice0' (Module coreir_slice)
  wire [15:0] slice0__in;
  wire [15:0] slice0__out;
  coreir_slice #(.hi(16),.lo(0),.width(16)) slice0(
    .in(slice0__in),
    .out(slice0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[15:0] = extendA__out[15:0];
  assign extendB__in[3:0] = B[3:0];
  assign op0__in1[15:0] = extendB__out[15:0];
  assign slice0__in[15:0] = op0__out[15:0];
  assign Y[15:0] = slice0__out[15:0];

endmodule //shr_U21

module __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__16 (
  input  cfg_clk,
  input [15:0] cfg_d,
  input  cfg_en,
  input  cfg_rst_n,
  input [15:0] data_in,
  output  debug_irq
);
  //Wire declarations for instance 'self__DOT__debug_irq__DOLLAR__bit_const_0' (Module corebit_const)
  wire  self__DOT__debug_irq__DOLLAR__bit_const_0__out;
  corebit_const #(.value(0)) self__DOT__debug_irq__DOLLAR__bit_const_0(
    .out(self__DOT__debug_irq__DOLLAR__bit_const_0__out)
  );

  //All the connections
  assign debug_irq = self__DOT__debug_irq__DOLLAR__bit_const_0__out;

endmodule //__DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__16

module coreir_neq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 != in1;

endmodule //coreir_neq

module __DOLLAR__paramod__BACKSLASH__test_lut__BACKSLASH__DataWidth__EQUALS__1 (
  input [7:0] cfg_a,
  input  cfg_clk,
  input [31:0] cfg_d,
  input  cfg_en,
  input  cfg_rst_n,
  input  op_a_in,
  input  op_b_in,
  input  op_c_in,
  output  res
);
  //All the connections
  assign res = op_a_in;

endmodule //__DOLLAR__paramod__BACKSLASH__test_lut__BACKSLASH__DataWidth__EQUALS__1

// module reg #(parameter clk_posedge=1, parameter init=1) (
//   input clk,
//   input in,
//   output out
// );
// reg outReg = init;
// always @(posedge clk) begin
//   outReg <= in;
// end
// assign out = outReg;

// endmodule //reg

module add_U2 (
  input [16:0] A,
  input [0:0] B,
  output [16:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [16:0] extendA__in;
  wire [16:0] extendA__out;
  coreir_zext #(.width_in(17),.width_out(17)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [16:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(17)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_add)
  wire [16:0] op0__in0;
  wire [16:0] op0__in1;
  wire [16:0] op0__out;
  coreir_add #(.width(17)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[16:0] = A[16:0];
  assign op0__in0[16:0] = extendA__out[16:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[16:0] = extendB__out[16:0];
  assign Y[16:0] = op0__out[16:0];

endmodule //add_U2

module __DOLLAR__paramod__BACKSLASH__test_full_add__BACKSLASH__DataWidth__EQUALS__16 (
  input [15:0] a,
  input [15:0] b,
  input  c_in,
  output  c_out,
  output [15:0] res
);
  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277' (Module add_U1)
  wire [15:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A;
  wire [15:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B;
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y;
  add_U1 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278' (Module add_U2)
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A;
  wire [0:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__B;
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y;
  add_U2 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y)
  );

  //All the connections
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__B[0] = c_in;
  assign c_out = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[16];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[0] = a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[1] = a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[10] = a[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[11] = a[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[12] = a[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[13] = a[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[14] = a[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[15] = a[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[2] = a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[3] = a[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[4] = a[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[5] = a[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[6] = a[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[7] = a[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[8] = a[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__A[9] = a[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[0] = b[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[1] = b[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[10] = b[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[11] = b[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[12] = b[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[13] = b[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[14] = b[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[15] = b[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[2] = b[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[3] = b[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[4] = b[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[5] = b[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[6] = b[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[7] = b[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[8] = b[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__B[9] = b[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[16];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__A[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__277__Y[9];
  assign res[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[0];
  assign res[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[1];
  assign res[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[10];
  assign res[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[11];
  assign res[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[12];
  assign res[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[13];
  assign res[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[14];
  assign res[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[15];
  assign res[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[2];
  assign res[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[3];
  assign res[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[4];
  assign res[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[5];
  assign res[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[6];
  assign res[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[7];
  assign res[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[8];
  assign res[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__278__Y[9];

endmodule //__DOLLAR__paramod__BACKSLASH__test_full_add__BACKSLASH__DataWidth__EQUALS__16

module test_full_add (
  input [15:0] a,
  input [15:0] b,
  input  c_in,
  output  c_out,
  output [15:0] res
);
  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33' (Module add_U1)
  wire [15:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A;
  wire [15:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B;
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y;
  add_U1 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34' (Module add_U2)
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A;
  wire [0:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__B;
  wire [16:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y;
  add_U2 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y)
  );

  //All the connections
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__B[0] = c_in;
  assign c_out = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[16];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[0] = a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[1] = a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[10] = a[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[11] = a[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[12] = a[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[13] = a[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[14] = a[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[15] = a[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[2] = a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[3] = a[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[4] = a[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[5] = a[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[6] = a[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[7] = a[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[8] = a[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__A[9] = a[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[0] = b[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[1] = b[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[10] = b[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[11] = b[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[12] = b[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[13] = b[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[14] = b[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[15] = b[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[2] = b[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[3] = b[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[4] = b[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[5] = b[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[6] = b[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[7] = b[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[8] = b[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__B[9] = b[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[10];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[11];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[12];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[13];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[14];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[15];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[16];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[3];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[4];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[5];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[6];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[7];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[8];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__A[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__33__Y[9];
  assign res[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[0];
  assign res[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[1];
  assign res[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[10];
  assign res[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[11];
  assign res[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[12];
  assign res[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[13];
  assign res[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[14];
  assign res[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[15];
  assign res[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[2];
  assign res[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[3];
  assign res[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[4];
  assign res[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[5];
  assign res[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[6];
  assign res[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[7];
  assign res[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[8];
  assign res[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_full_add__DOT__sv__COLON__50__DOLLAR__34__Y[9];

endmodule //test_full_add

module reg_arst #(parameter arst_posedge=1, parameter clk_posedge=1, parameter init=1) (
  input clk,
  input in,
  input arst,
  output out
);
reg outReg;
wire real_rst;
assign real_rst = arst_posedge ? arst : ~arst;
wire real_clk;
assign real_clk = clk_posedge ? clk : ~clk;
always @(posedge real_clk, posedge real_rst) begin
  if (real_rst) outReg <= init;
  else outReg <= in;
end
assign out = outReg;

endmodule //reg_arst

module reduce_and_U44 (
  input [7:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_andr)
  wire [7:0] op0__in;
  wire  op0__out;
  coreir_andr #(.width(8)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[7:0] = A[7:0];
  assign Y[0] = op0__out;

endmodule //reduce_and_U44

module adff_U24 #(parameter init=1) (
  input  ARST,
  input  CLK,
  input [15:0] D,
  output [15:0] Q
);
  //Wire declarations for instance 'reg0' (Module coreir_reg_arst)
  wire  reg0__arst;
  wire  reg0__clk;
  wire [15:0] reg0__in;
  wire [15:0] reg0__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(init),.width(16)) reg0(
    .arst(reg0__arst),
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //Wire declarations for instance 'toClk0' (Module coreir_wrap)
  wire  toClk0__in;
  wire  toClk0__out;
  coreir_wrap toClk0(
    .in(toClk0__in),
    .out(toClk0__out)
  );

  //Wire declarations for instance 'toRST0' (Module coreir_wrap)
  wire  toRST0__in;
  wire  toRST0__out;
  coreir_wrap toRST0(
    .in(toRST0__in),
    .out(toRST0__out)
  );

  //All the connections
  assign reg0__arst = toRST0__out;
  assign reg0__clk = toClk0__out;
  assign reg0__in[15:0] = D[15:0];
  assign Q[15:0] = reg0__out[15:0];
  assign toRST0__in = ARST;
  assign toClk0__in = CLK;

endmodule //adff_U24

module adff_U25 #(parameter init=1) (
  input  ARST,
  input  CLK,
  input [63:0] D,
  output [63:0] Q
);
  //Wire declarations for instance 'reg0' (Module coreir_reg_arst)
  wire  reg0__arst;
  wire  reg0__clk;
  wire [63:0] reg0__in;
  wire [63:0] reg0__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(init),.width(64)) reg0(
    .arst(reg0__arst),
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //Wire declarations for instance 'toClk0' (Module coreir_wrap)
  wire  toClk0__in;
  wire  toClk0__out;
  coreir_wrap toClk0(
    .in(toClk0__in),
    .out(toClk0__out)
  );

  //Wire declarations for instance 'toRST0' (Module coreir_wrap)
  wire  toRST0__in;
  wire  toRST0__out;
  coreir_wrap toRST0(
    .in(toRST0__in),
    .out(toRST0__out)
  );

  //All the connections
  assign reg0__arst = toRST0__out;
  assign reg0__clk = toClk0__out;
  assign reg0__in[63:0] = D[63:0];
  assign Q[63:0] = reg0__out[63:0];
  assign toRST0__in = ARST;
  assign toClk0__in = CLK;

endmodule //adff_U25

module adff_U7 #(parameter init=1) (
  input  ARST,
  input  CLK,
  input [0:0] D,
  output [0:0] Q
);
  //Wire declarations for instance 'reg0' (Module coreir_reg_arst)
  wire  reg0__arst;
  wire  reg0__clk;
  wire [0:0] reg0__in;
  wire [0:0] reg0__out;
  coreir_reg_arst #(.arst_posedge(0),.clk_posedge(1),.init(init),.width(1)) reg0(
    .arst(reg0__arst),
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //Wire declarations for instance 'toClk0' (Module coreir_wrap)
  wire  toClk0__in;
  wire  toClk0__out;
  coreir_wrap toClk0(
    .in(toClk0__in),
    .out(toClk0__out)
  );

  //Wire declarations for instance 'toRST0' (Module coreir_wrap)
  wire  toRST0__in;
  wire  toRST0__out;
  coreir_wrap toRST0(
    .in(toRST0__in),
    .out(toRST0__out)
  );

  //All the connections
  assign reg0__arst = toRST0__out;
  assign reg0__clk = toClk0__out;
  assign reg0__in[0:0] = D[0:0];
  assign Q[0:0] = reg0__out[0:0];
  assign toRST0__in = ARST;
  assign toClk0__in = CLK;

endmodule //adff_U7

module adff_U9 #(parameter init=1) (
  input  ARST,
  input  CLK,
  input [15:0] D,
  output [15:0] Q
);
  //Wire declarations for instance 'reg0' (Module coreir_reg_arst)
  wire  reg0__arst;
  wire  reg0__clk;
  wire [15:0] reg0__in;
  wire [15:0] reg0__out;
  coreir_reg_arst #(.arst_posedge(0),.clk_posedge(1),.init(init),.width(16)) reg0(
    .arst(reg0__arst),
    .clk(reg0__clk),
    .in(reg0__in),
    .out(reg0__out)
  );

  //Wire declarations for instance 'toClk0' (Module coreir_wrap)
  wire  toClk0__in;
  wire  toClk0__out;
  coreir_wrap toClk0(
    .in(toClk0__in),
    .out(toClk0__out)
  );

  //Wire declarations for instance 'toRST0' (Module coreir_wrap)
  wire  toRST0__in;
  wire  toRST0__out;
  coreir_wrap toRST0(
    .in(toRST0__in),
    .out(toRST0__out)
  );

  //All the connections
  assign reg0__arst = toRST0__out;
  assign reg0__clk = toClk0__out;
  assign reg0__in[15:0] = D[15:0];
  assign Q[15:0] = reg0__out[15:0];
  assign toRST0__in = ARST;
  assign toClk0__in = CLK;

endmodule //adff_U9

module xor_U27 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_xor)
  wire [0:0] op0__in0;
  wire [0:0] op0__in1;
  wire [0:0] op0__out;
  coreir_xor #(.width(1)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in0[0:0] = extendA__out[0:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[0:0] = extendB__out[0:0];
  assign Y[0:0] = op0__out[0:0];

endmodule //xor_U27

module and_U28 (
  input [15:0] A,
  input [15:0] B,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [15:0] extendB__in;
  wire [15:0] extendB__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_and)
  wire [15:0] op0__in0;
  wire [15:0] op0__in1;
  wire [15:0] op0__out;
  coreir_and #(.width(16)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[15:0] = extendA__out[15:0];
  assign extendB__in[15:0] = B[15:0];
  assign op0__in1[15:0] = extendB__out[15:0];
  assign Y[15:0] = op0__out[15:0];

endmodule //and_U28

module and_U3 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_and)
  wire [0:0] op0__in0;
  wire [0:0] op0__in1;
  wire [0:0] op0__out;
  coreir_and #(.width(1)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in0[0:0] = extendA__out[0:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[0:0] = extendB__out[0:0];
  assign Y[0:0] = op0__out[0:0];

endmodule //and_U3

module test_mult_add (
  input [15:0] a,
  input [15:0] b,
  output  c_out,
  input  is_signed,
  output [31:0] res
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__Y)
  );

  //Wire declarations for instance '__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37' (Module mul_U4)
  wire [16:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A;
  wire [16:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B;
  wire [33:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y;
  mul_U4 __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37(
    .A(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A),
    .B(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B),
    .Y(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y)
  );

  //Wire declarations for instance 'self__DOT__c_out__DOLLAR__bit_const_0' (Module corebit_const)
  wire  self__DOT__c_out__DOLLAR__bit_const_0__out;
  corebit_const #(.value(0)) self__DOT__c_out__DOLLAR__bit_const_0(
    .out(self__DOT__c_out__DOLLAR__bit_const_0__out)
  );

  //All the connections
  assign c_out = self__DOT__c_out__DOLLAR__bit_const_0__out;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__A[0] = is_signed;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__A[0] = is_signed;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__B[0] = a[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[16] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__35__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__B[0] = b[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[16] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__36__Y[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[0] = a[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[1] = a[1];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[10] = a[10];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[11] = a[11];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[12] = a[12];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[13] = a[13];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[14] = a[14];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[15] = a[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[2] = a[2];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[3] = a[3];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[4] = a[4];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[5] = a[5];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[6] = a[6];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[7] = a[7];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[8] = a[8];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__A[9] = a[9];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[0] = b[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[1] = b[1];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[10] = b[10];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[11] = b[11];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[12] = b[12];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[13] = b[13];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[14] = b[14];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[15] = b[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[2] = b[2];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[3] = b[3];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[4] = b[4];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[5] = b[5];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[6] = b[6];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[7] = b[7];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[8] = b[8];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__B[9] = b[9];
  assign res[0] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[0];
  assign res[1] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[1];
  assign res[10] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[10];
  assign res[11] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[11];
  assign res[12] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[12];
  assign res[13] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[13];
  assign res[14] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[14];
  assign res[15] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[15];
  assign res[16] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[16];
  assign res[17] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[17];
  assign res[18] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[18];
  assign res[19] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[19];
  assign res[2] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[2];
  assign res[20] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[20];
  assign res[21] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[21];
  assign res[22] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[22];
  assign res[23] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[23];
  assign res[24] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[24];
  assign res[25] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[25];
  assign res[26] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[26];
  assign res[27] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[27];
  assign res[28] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[28];
  assign res[29] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[29];
  assign res[3] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[3];
  assign res[30] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[30];
  assign res[31] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[31];
  assign res[4] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[4];
  assign res[5] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[5];
  assign res[6] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[6];
  assign res[7] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[7];
  assign res[8] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[8];
  assign res[9] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__37__Y[9];

endmodule //test_mult_add

module __DOLLAR__paramod__BACKSLASH__test_mult_add__BACKSLASH__DataWidth__EQUALS__16 (
  input [15:0] a,
  input [15:0] b,
  output  c_out,
  input  is_signed,
  output [31:0] res
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__Y)
  );

  //Wire declarations for instance '__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286' (Module mul_U4)
  wire [16:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A;
  wire [16:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B;
  wire [33:0] __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y;
  mul_U4 __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286(
    .A(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A),
    .B(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B),
    .Y(__DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y)
  );

  //Wire declarations for instance 'self__DOT__c_out__DOLLAR__bit_const_0' (Module corebit_const)
  wire  self__DOT__c_out__DOLLAR__bit_const_0__out;
  corebit_const #(.value(0)) self__DOT__c_out__DOLLAR__bit_const_0(
    .out(self__DOT__c_out__DOLLAR__bit_const_0__out)
  );

  //All the connections
  assign c_out = self__DOT__c_out__DOLLAR__bit_const_0__out;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__A[0] = is_signed;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__A[0] = is_signed;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__B[0] = a[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[16] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__61__DOLLAR__284__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__B[0] = b[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[16] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__62__DOLLAR__285__Y[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[0] = a[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[1] = a[1];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[10] = a[10];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[11] = a[11];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[12] = a[12];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[13] = a[13];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[14] = a[14];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[15] = a[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[2] = a[2];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[3] = a[3];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[4] = a[4];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[5] = a[5];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[6] = a[6];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[7] = a[7];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[8] = a[8];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__A[9] = a[9];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[0] = b[0];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[1] = b[1];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[10] = b[10];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[11] = b[11];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[12] = b[12];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[13] = b[13];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[14] = b[14];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[15] = b[15];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[2] = b[2];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[3] = b[3];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[4] = b[4];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[5] = b[5];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[6] = b[6];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[7] = b[7];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[8] = b[8];
  assign __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__B[9] = b[9];
  assign res[0] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[0];
  assign res[1] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[1];
  assign res[10] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[10];
  assign res[11] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[11];
  assign res[12] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[12];
  assign res[13] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[13];
  assign res[14] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[14];
  assign res[15] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[15];
  assign res[16] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[16];
  assign res[17] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[17];
  assign res[18] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[18];
  assign res[19] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[19];
  assign res[2] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[2];
  assign res[20] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[20];
  assign res[21] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[21];
  assign res[22] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[22];
  assign res[23] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[23];
  assign res[24] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[24];
  assign res[25] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[25];
  assign res[26] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[26];
  assign res[27] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[27];
  assign res[28] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[28];
  assign res[29] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[29];
  assign res[3] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[3];
  assign res[30] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[30];
  assign res[31] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[31];
  assign res[4] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[4];
  assign res[5] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[5];
  assign res[6] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[6];
  assign res[7] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[7];
  assign res[8] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[8];
  assign res[9] = __DOLLAR__mul__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_mult_add__DOT__sv__COLON__64__DOLLAR__286__Y[9];

endmodule //__DOLLAR__paramod__BACKSLASH__test_mult_add__BACKSLASH__DataWidth__EQUALS__16

module and_U42 (
  input [1:0] A,
  input [1:0] B,
  output [1:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [1:0] extendA__in;
  wire [1:0] extendA__out;
  coreir_zext #(.width_in(2),.width_out(2)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [1:0] extendB__in;
  wire [1:0] extendB__out;
  coreir_zext #(.width_in(2),.width_out(2)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_and)
  wire [1:0] op0__in0;
  wire [1:0] op0__in1;
  wire [1:0] op0__out;
  coreir_and #(.width(2)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[1:0] = A[1:0];
  assign op0__in0[1:0] = extendA__out[1:0];
  assign extendB__in[1:0] = B[1:0];
  assign op0__in1[1:0] = extendB__out[1:0];
  assign Y[1:0] = op0__out[1:0];

endmodule //and_U42

module eq_U15 (
  input [3:0] A,
  input [3:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [3:0] extendA__in;
  wire [3:0] extendA__out;
  coreir_zext #(.width_in(4),.width_out(4)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [3:0] extendB__in;
  wire [3:0] extendB__out;
  coreir_zext #(.width_in(4),.width_out(4)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [3:0] op0__in0;
  wire [3:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(4)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[3:0] = A[3:0];
  assign op0__in0[3:0] = extendA__out[3:0];
  assign extendB__in[3:0] = B[3:0];
  assign op0__in1[3:0] = extendB__out[3:0];
  assign Y[0] = op0__out;

endmodule //eq_U15

module rtMux_U26 (
  input [31:0] A,
  input [31:0] B,
  input  S,
  output [31:0] Y
);
  //Wire declarations for instance 'mux0' (Module coreir_mux)
  wire [31:0] mux0__in0;
  wire [31:0] mux0__in1;
  wire [31:0] mux0__out;
  wire  mux0__sel;
  coreir_mux #(.width(32)) mux0(
    .in0(mux0__in0),
    .in1(mux0__in1),
    .out(mux0__out),
    .sel(mux0__sel)
  );

  //All the connections
  assign mux0__in0[31:0] = A[31:0];
  assign mux0__in1[31:0] = B[31:0];
  assign Y[31:0] = mux0__out[31:0];
  assign mux0__sel = S;

endmodule //rtMux_U26

module eq_U16 (
  input [31:0] A,
  input [31:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [31:0] extendA__in;
  wire [31:0] extendA__out;
  coreir_zext #(.width_in(32),.width_out(32)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [31:0] extendB__in;
  wire [31:0] extendB__out;
  coreir_zext #(.width_in(32),.width_out(32)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [31:0] op0__in0;
  wire [31:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(32)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[31:0] = A[31:0];
  assign op0__in0[31:0] = extendA__out[31:0];
  assign extendB__in[31:0] = B[31:0];
  assign op0__in1[31:0] = extendB__out[31:0];
  assign Y[0] = op0__out;

endmodule //eq_U16

module eq_U23 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [0:0] op0__in0;
  wire [0:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(1)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in0[0:0] = extendA__out[0:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[0:0] = extendB__out[0:0];
  assign Y[0] = op0__out;

endmodule //eq_U23

module eq_U5 (
  input [1:0] A,
  input [1:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [1:0] extendA__in;
  wire [1:0] extendA__out;
  coreir_zext #(.width_in(2),.width_out(2)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [1:0] extendB__in;
  wire [1:0] extendB__out;
  coreir_zext #(.width_in(2),.width_out(2)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_eq)
  wire [1:0] op0__in0;
  wire [1:0] op0__in1;
  wire  op0__out;
  coreir_eq #(.width(2)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[1:0] = A[1:0];
  assign op0__in0[1:0] = extendA__out[1:0];
  assign extendB__in[1:0] = B[1:0];
  assign op0__in1[1:0] = extendB__out[1:0];
  assign Y[0] = op0__out;

endmodule //eq_U5

module logic_and_U19 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'aRed' (Module coreir_orr)
  wire [0:0] aRed__in;
  wire  aRed__out;
  coreir_orr #(.width(1)) aRed(
    .in(aRed__in),
    .out(aRed__out)
  );

  //Wire declarations for instance 'andOps' (Module corebit_and)
  wire  andOps__in0;
  wire  andOps__in1;
  wire  andOps__out;
  corebit_and andOps(
    .in0(andOps__in0),
    .in1(andOps__in1),
    .out(andOps__out)
  );

  //Wire declarations for instance 'bRed' (Module coreir_orr)
  wire [0:0] bRed__in;
  wire  bRed__out;
  coreir_orr #(.width(1)) bRed(
    .in(bRed__in),
    .out(bRed__out)
  );

  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //All the connections
  assign aRed__in[0:0] = extendA__out[0:0];
  assign andOps__in0 = aRed__out;
  assign andOps__in1 = bRed__out;
  assign Y[0] = andOps__out;
  assign bRed__in[0:0] = extendB__out[0:0];
  assign extendA__in[0:0] = A[0:0];
  assign extendB__in[0:0] = B[0:0];

endmodule //logic_and_U19

module logic_not_U33 (
  input [0:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'negate' (Module corebit_not)
  wire  negate__in;
  wire  negate__out;
  corebit_not negate(
    .in(negate__in),
    .out(negate__out)
  );

  //Wire declarations for instance 'reduce' (Module coreir_orr)
  wire [0:0] reduce__in;
  wire  reduce__out;
  coreir_orr #(.width(1)) reduce(
    .in(reduce__in),
    .out(reduce__out)
  );

  //All the connections
  assign negate__in = reduce__out;
  assign Y[0] = negate__out;
  assign reduce__in[0:0] = A[0:0];

endmodule //logic_not_U33

module ne_U34 (
  input [0:0] A,
  input [0:0] B,
  output [0:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [0:0] extendA__in;
  wire [0:0] extendA__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [0:0] extendB__in;
  wire [0:0] extendB__out;
  coreir_zext #(.width_in(1),.width_out(1)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_neq)
  wire [0:0] op0__in0;
  wire [0:0] op0__in1;
  wire  op0__out;
  coreir_neq #(.width(1)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[0:0] = A[0:0];
  assign op0__in0[0:0] = extendA__out[0:0];
  assign extendB__in[0:0] = B[0:0];
  assign op0__in1[0:0] = extendB__out[0:0];
  assign Y[0] = op0__out;

endmodule //ne_U34

module or_U36 (
  input [15:0] A,
  input [15:0] B,
  output [15:0] Y
);
  //Wire declarations for instance 'extendA' (Module coreir_zext)
  wire [15:0] extendA__in;
  wire [15:0] extendA__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendA(
    .in(extendA__in),
    .out(extendA__out)
  );

  //Wire declarations for instance 'extendB' (Module coreir_zext)
  wire [15:0] extendB__in;
  wire [15:0] extendB__out;
  coreir_zext #(.width_in(16),.width_out(16)) extendB(
    .in(extendB__in),
    .out(extendB__out)
  );

  //Wire declarations for instance 'op0' (Module coreir_or)
  wire [15:0] op0__in0;
  wire [15:0] op0__in1;
  wire [15:0] op0__out;
  coreir_or #(.width(16)) op0(
    .in0(op0__in0),
    .in1(op0__in1),
    .out(op0__out)
  );

  //All the connections
  assign extendA__in[15:0] = A[15:0];
  assign op0__in0[15:0] = extendA__out[15:0];
  assign extendB__in[15:0] = B[15:0];
  assign op0__in1[15:0] = extendB__out[15:0];
  assign Y[15:0] = op0__out[15:0];

endmodule //or_U36

module reduce_or_U12 (
  input [2:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [2:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(3)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[2:0] = A[2:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U12

module reduce_or_U13 (
  input [1:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [1:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(2)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[1:0] = A[1:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U13

module reduce_or_U31 (
  input [14:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [14:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(15)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[14:0] = A[14:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U31

module reduce_or_U38 (
  input [0:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [0:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(1)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[0:0] = A[0:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U38

module reduce_or_U39 (
  input [31:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [31:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(32)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[31:0] = A[31:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U39

module reduce_or_U43 (
  input [9:0] A,
  output [0:0] Y
);
  //Wire declarations for instance 'op0' (Module coreir_orr)
  wire [9:0] op0__in;
  wire  op0__out;
  coreir_orr #(.width(10)) op0(
    .in(op0__in),
    .out(op0__out)
  );

  //All the connections
  assign op0__in[9:0] = A[9:0];
  assign Y[0] = op0__out;

endmodule //reduce_or_U43

module rtMux_U10 (
  input [15:0] A,
  input [15:0] B,
  input  S,
  output [15:0] Y
);
  //Wire declarations for instance 'mux0' (Module coreir_mux)
  wire [15:0] mux0__in0;
  wire [15:0] mux0__in1;
  wire [15:0] mux0__out;
  wire  mux0__sel;
  coreir_mux #(.width(16)) mux0(
    .in0(mux0__in0),
    .in1(mux0__in1),
    .out(mux0__out),
    .sel(mux0__sel)
  );

  //All the connections
  assign mux0__in0[15:0] = A[15:0];
  assign mux0__in1[15:0] = B[15:0];
  assign Y[15:0] = mux0__out[15:0];
  assign mux0__sel = S;

endmodule //rtMux_U10

module sb_unq1 (
  input  clk,
  input [31:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  output [63:0] config_sb_res,
  input [15:0] in_0_0,
  input [15:0] in_0_1,
  input [15:0] in_0_2,
  input [15:0] in_0_3,
  input [15:0] in_0_4,
  input [15:0] in_1_0,
  input [15:0] in_1_1,
  input [15:0] in_1_2,
  input [15:0] in_1_3,
  input [15:0] in_1_4,
  input [15:0] in_2_0,
  input [15:0] in_2_1,
  input [15:0] in_2_2,
  input [15:0] in_2_3,
  input [15:0] in_2_4,
  input [15:0] in_3_0,
  input [15:0] in_3_1,
  input [15:0] in_3_2,
  input [15:0] in_3_3,
  input [15:0] in_3_4,
  output [15:0] out_0_0,
  output [15:0] out_0_1,
  output [15:0] out_0_2,
  output [15:0] out_0_3,
  output [15:0] out_0_4,
  output [15:0] out_1_0,
  output [15:0] out_1_1,
  output [15:0] out_1_2,
  output [15:0] out_1_3,
  output [15:0] out_1_4,
  output [15:0] out_2_0,
  output [15:0] out_2_1,
  output [15:0] out_2_2,
  output [15:0] out_2_3,
  output [15:0] out_2_4,
  output [15:0] out_3_0,
  output [15:0] out_3_1,
  output [15:0] out_3_2,
  output [15:0] out_3_3,
  output [15:0] out_3_4,
  input [15:0] pe_output_0,
  input  reset
);
  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196(
    .A(__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__731' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__731__ARST;
  wire  __DOLLAR__procdff__DOLLAR__731__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__731__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__731__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__731(
    .ARST(__DOLLAR__procdff__DOLLAR__731__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__731__CLK),
    .D(__DOLLAR__procdff__DOLLAR__731__D),
    .Q(__DOLLAR__procdff__DOLLAR__731__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__732' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__732__ARST;
  wire  __DOLLAR__procdff__DOLLAR__732__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__732__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__732__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__732(
    .ARST(__DOLLAR__procdff__DOLLAR__732__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__732__CLK),
    .D(__DOLLAR__procdff__DOLLAR__732__D),
    .Q(__DOLLAR__procdff__DOLLAR__732__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__733' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__733__ARST;
  wire  __DOLLAR__procdff__DOLLAR__733__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__733__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__733__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__733(
    .ARST(__DOLLAR__procdff__DOLLAR__733__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__733__CLK),
    .D(__DOLLAR__procdff__DOLLAR__733__D),
    .Q(__DOLLAR__procdff__DOLLAR__733__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__734' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__734__ARST;
  wire  __DOLLAR__procdff__DOLLAR__734__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__734__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__734__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__734(
    .ARST(__DOLLAR__procdff__DOLLAR__734__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__734__CLK),
    .D(__DOLLAR__procdff__DOLLAR__734__D),
    .Q(__DOLLAR__procdff__DOLLAR__734__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__735' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__735__ARST;
  wire  __DOLLAR__procdff__DOLLAR__735__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__735__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__735__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__735(
    .ARST(__DOLLAR__procdff__DOLLAR__735__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__735__CLK),
    .D(__DOLLAR__procdff__DOLLAR__735__D),
    .Q(__DOLLAR__procdff__DOLLAR__735__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__736' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__736__ARST;
  wire  __DOLLAR__procdff__DOLLAR__736__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__736__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__736__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__736(
    .ARST(__DOLLAR__procdff__DOLLAR__736__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__736__CLK),
    .D(__DOLLAR__procdff__DOLLAR__736__D),
    .Q(__DOLLAR__procdff__DOLLAR__736__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__737' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__737__ARST;
  wire  __DOLLAR__procdff__DOLLAR__737__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__737__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__737__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__737(
    .ARST(__DOLLAR__procdff__DOLLAR__737__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__737__CLK),
    .D(__DOLLAR__procdff__DOLLAR__737__D),
    .Q(__DOLLAR__procdff__DOLLAR__737__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__738' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__738__ARST;
  wire  __DOLLAR__procdff__DOLLAR__738__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__738__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__738__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__738(
    .ARST(__DOLLAR__procdff__DOLLAR__738__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__738__CLK),
    .D(__DOLLAR__procdff__DOLLAR__738__D),
    .Q(__DOLLAR__procdff__DOLLAR__738__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__739' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__739__ARST;
  wire  __DOLLAR__procdff__DOLLAR__739__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__739__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__739__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__739(
    .ARST(__DOLLAR__procdff__DOLLAR__739__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__739__CLK),
    .D(__DOLLAR__procdff__DOLLAR__739__D),
    .Q(__DOLLAR__procdff__DOLLAR__739__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__740' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__740__ARST;
  wire  __DOLLAR__procdff__DOLLAR__740__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__740__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__740__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__740(
    .ARST(__DOLLAR__procdff__DOLLAR__740__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__740__CLK),
    .D(__DOLLAR__procdff__DOLLAR__740__D),
    .Q(__DOLLAR__procdff__DOLLAR__740__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__741' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__741__ARST;
  wire  __DOLLAR__procdff__DOLLAR__741__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__741__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__741__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__741(
    .ARST(__DOLLAR__procdff__DOLLAR__741__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__741__CLK),
    .D(__DOLLAR__procdff__DOLLAR__741__D),
    .Q(__DOLLAR__procdff__DOLLAR__741__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__742' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__742__ARST;
  wire  __DOLLAR__procdff__DOLLAR__742__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__742__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__742__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__742(
    .ARST(__DOLLAR__procdff__DOLLAR__742__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__742__CLK),
    .D(__DOLLAR__procdff__DOLLAR__742__D),
    .Q(__DOLLAR__procdff__DOLLAR__742__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__743' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__743__ARST;
  wire  __DOLLAR__procdff__DOLLAR__743__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__743__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__743__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__743(
    .ARST(__DOLLAR__procdff__DOLLAR__743__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__743__CLK),
    .D(__DOLLAR__procdff__DOLLAR__743__D),
    .Q(__DOLLAR__procdff__DOLLAR__743__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__744' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__744__ARST;
  wire  __DOLLAR__procdff__DOLLAR__744__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__744__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__744__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__744(
    .ARST(__DOLLAR__procdff__DOLLAR__744__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__744__CLK),
    .D(__DOLLAR__procdff__DOLLAR__744__D),
    .Q(__DOLLAR__procdff__DOLLAR__744__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__745' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__745__ARST;
  wire  __DOLLAR__procdff__DOLLAR__745__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__745__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__745__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__745(
    .ARST(__DOLLAR__procdff__DOLLAR__745__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__745__CLK),
    .D(__DOLLAR__procdff__DOLLAR__745__D),
    .Q(__DOLLAR__procdff__DOLLAR__745__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__746' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__746__ARST;
  wire  __DOLLAR__procdff__DOLLAR__746__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__746__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__746__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__746(
    .ARST(__DOLLAR__procdff__DOLLAR__746__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__746__CLK),
    .D(__DOLLAR__procdff__DOLLAR__746__D),
    .Q(__DOLLAR__procdff__DOLLAR__746__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__747' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__747__ARST;
  wire  __DOLLAR__procdff__DOLLAR__747__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__747__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__747__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__747(
    .ARST(__DOLLAR__procdff__DOLLAR__747__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__747__CLK),
    .D(__DOLLAR__procdff__DOLLAR__747__D),
    .Q(__DOLLAR__procdff__DOLLAR__747__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__748' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__748__ARST;
  wire  __DOLLAR__procdff__DOLLAR__748__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__748__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__748__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__748(
    .ARST(__DOLLAR__procdff__DOLLAR__748__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__748__CLK),
    .D(__DOLLAR__procdff__DOLLAR__748__D),
    .Q(__DOLLAR__procdff__DOLLAR__748__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__749' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__749__ARST;
  wire  __DOLLAR__procdff__DOLLAR__749__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__749__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__749__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__749(
    .ARST(__DOLLAR__procdff__DOLLAR__749__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__749__CLK),
    .D(__DOLLAR__procdff__DOLLAR__749__D),
    .Q(__DOLLAR__procdff__DOLLAR__749__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__750' (Module adff_U24)
  wire  __DOLLAR__procdff__DOLLAR__750__ARST;
  wire  __DOLLAR__procdff__DOLLAR__750__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__750__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__750__Q;
  adff_U24 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__750(
    .ARST(__DOLLAR__procdff__DOLLAR__750__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__750__CLK),
    .D(__DOLLAR__procdff__DOLLAR__750__D),
    .Q(__DOLLAR__procdff__DOLLAR__750__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__751' (Module adff_U25)
  wire  __DOLLAR__procdff__DOLLAR__751__ARST;
  wire  __DOLLAR__procdff__DOLLAR__751__CLK;
  wire [63:0] __DOLLAR__procdff__DOLLAR__751__D;
  wire [63:0] __DOLLAR__procdff__DOLLAR__751__Q;
  adff_U25 #(.init(64'b0000000000000000000000001111111111111111111111111111111111111111)) __DOLLAR__procdff__DOLLAR__751(
    .ARST(__DOLLAR__procdff__DOLLAR__751__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__751__CLK),
    .D(__DOLLAR__procdff__DOLLAR__751__D),
    .Q(__DOLLAR__procdff__DOLLAR__751__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__412_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__412_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__412_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__412_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__412_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__412_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__412_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__412_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__413_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__413_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__413_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__413_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__413_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__413_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__413_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__413_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__414_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__414_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__414_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__414_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__414_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__414_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__414_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__414_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__415_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__415_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__415_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__415_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__415_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__415_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__415_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__415_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__417_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__417_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__417_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__417_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__417_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__417_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__417_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__417_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__418_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__418_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__418_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__418_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__418_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__418_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__418_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__418_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__419_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__419_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__419_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__419_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__419_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__419_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__419_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__419_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__420_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__420_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__420_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__420_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__420_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__420_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__420_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__420_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__422_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__422_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__422_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__422_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__422_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__422_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__422_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__422_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__423_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__423_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__423_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__423_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__423_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__423_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__423_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__423_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__424_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__424_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__424_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__424_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__424_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__424_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__424_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__424_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__425_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__425_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__425_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__425_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__425_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__425_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__425_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__425_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__427_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__427_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__427_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__427_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__427_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__427_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__427_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__427_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__428_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__428_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__428_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__428_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__428_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__428_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__428_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__428_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__429_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__429_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__429_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__429_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__429_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__429_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__429_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__429_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__430_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__430_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__430_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__430_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__430_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__430_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__430_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__430_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__432_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__432_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__432_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__432_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__432_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__432_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__432_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__432_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__433_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__433_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__433_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__433_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__433_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__433_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__433_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__433_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__434_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__434_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__434_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__434_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__434_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__434_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__434_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__434_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__435_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__435_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__435_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__435_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__435_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__435_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__435_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__435_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__437_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__437_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__437_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__437_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__437_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__437_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__437_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__437_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__438_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__438_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__438_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__438_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__438_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__438_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__438_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__438_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__439_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__439_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__439_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__439_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__439_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__439_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__439_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__439_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__440_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__440_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__440_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__440_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__440_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__440_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__440_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__440_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__442_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__442_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__442_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__442_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__442_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__442_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__442_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__442_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__443_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__443_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__443_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__443_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__443_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__443_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__443_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__443_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__444_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__444_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__444_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__444_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__444_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__444_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__444_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__444_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__445_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__445_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__445_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__445_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__445_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__445_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__445_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__445_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__447_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__447_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__447_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__447_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__447_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__447_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__447_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__447_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__448_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__448_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__448_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__448_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__448_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__448_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__448_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__448_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__449_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__449_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__449_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__449_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__449_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__449_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__449_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__449_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__450_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__450_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__450_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__450_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__450_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__450_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__450_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__450_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__452_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__452_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__452_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__452_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__452_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__452_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__452_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__452_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__453_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__453_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__453_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__453_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__453_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__453_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__453_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__453_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__454_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__454_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__454_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__454_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__454_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__454_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__454_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__454_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__455_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__455_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__455_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__455_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__455_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__455_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__455_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__455_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__457_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__457_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__457_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__457_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__457_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__457_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__457_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__457_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__458_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__458_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__458_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__458_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__458_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__458_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__458_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__458_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__459_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__459_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__459_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__459_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__459_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__459_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__459_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__459_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__460_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__460_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__460_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__460_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__460_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__460_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__460_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__460_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__462_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__462_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__462_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__462_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__462_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__462_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__462_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__462_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__463_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__463_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__463_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__463_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__463_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__463_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__463_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__463_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__464_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__464_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__464_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__464_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__464_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__464_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__464_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__464_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__465_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__465_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__465_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__465_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__465_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__465_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__465_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__465_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__467_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__467_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__467_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__467_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__467_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__467_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__467_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__467_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__468_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__468_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__468_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__468_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__468_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__468_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__468_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__468_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__469_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__469_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__469_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__469_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__469_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__469_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__469_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__469_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__470_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__470_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__470_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__470_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__470_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__470_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__470_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__470_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__472_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__472_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__472_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__472_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__472_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__472_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__472_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__472_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__473_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__473_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__473_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__473_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__473_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__473_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__473_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__473_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__474_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__474_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__474_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__474_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__474_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__474_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__474_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__474_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__475_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__475_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__475_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__475_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__475_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__475_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__475_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__475_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__477_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__477_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__477_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__477_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__477_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__477_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__477_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__477_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__478_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__478_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__478_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__478_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__478_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__478_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__478_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__478_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__479_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__479_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__479_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__479_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__479_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__479_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__479_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__479_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__480_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__480_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__480_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__480_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__480_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__480_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__480_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__480_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__482_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__482_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__482_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__482_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__482_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__482_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__482_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__482_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__483_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__483_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__483_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__483_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__483_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__483_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__483_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__483_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__484_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__484_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__484_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__484_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__484_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__484_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__484_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__484_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__485_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__485_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__485_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__485_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__485_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__485_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__485_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__485_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__487_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__487_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__487_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__487_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__487_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__487_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__487_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__487_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__488_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__488_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__488_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__488_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__488_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__488_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__488_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__488_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__489_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__489_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__489_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__489_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__489_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__489_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__489_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__489_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__490_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__490_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__490_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__490_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__490_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__490_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__490_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__490_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__492_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__492_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__492_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__492_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__492_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__492_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__492_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__492_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__493_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__493_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__493_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__493_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__493_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__493_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__493_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__493_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__494_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__494_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__494_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__494_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__494_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__494_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__494_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__494_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__495_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__495_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__495_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__495_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__495_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__495_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__495_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__495_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__497_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__497_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__497_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__497_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__497_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__497_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__497_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__497_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__498_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__498_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__498_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__498_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__498_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__498_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__498_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__498_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__499_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__499_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__499_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__499_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__499_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__499_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__499_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__499_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__500_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__500_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__500_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__500_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__500_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__500_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__500_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__500_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__502_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__502_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__502_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__502_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__502_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__502_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__502_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__502_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__503_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__503_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__503_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__503_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__503_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__503_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__503_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__503_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__504_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__504_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__504_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__504_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__504_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__504_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__504_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__504_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__505_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__505_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__505_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__505_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__505_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__505_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__505_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__505_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__507_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__507_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__507_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__507_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__507_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__507_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__507_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__507_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__508_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__508_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__508_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__508_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__508_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__508_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__508_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__508_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__509_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__509_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__509_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__509_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__509_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__509_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__509_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__509_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__510_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__510_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__510_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__510_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__510_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__510_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__510_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__510_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__513' (Module rtMux_U26)
  wire [31:0] __DOLLAR__procmux__DOLLAR__513__A;
  wire [31:0] __DOLLAR__procmux__DOLLAR__513__B;
  wire  __DOLLAR__procmux__DOLLAR__513__S;
  wire [31:0] __DOLLAR__procmux__DOLLAR__513__Y;
  rtMux_U26 __DOLLAR__procmux__DOLLAR__513(
    .A(__DOLLAR__procmux__DOLLAR__513__A),
    .B(__DOLLAR__procmux__DOLLAR__513__B),
    .S(__DOLLAR__procmux__DOLLAR__513__S),
    .Y(__DOLLAR__procmux__DOLLAR__513__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__514_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__514_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__514_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__514_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__514_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__514_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__514_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__515' (Module rtMux_U26)
  wire [31:0] __DOLLAR__procmux__DOLLAR__515__A;
  wire [31:0] __DOLLAR__procmux__DOLLAR__515__B;
  wire  __DOLLAR__procmux__DOLLAR__515__S;
  wire [31:0] __DOLLAR__procmux__DOLLAR__515__Y;
  rtMux_U26 __DOLLAR__procmux__DOLLAR__515(
    .A(__DOLLAR__procmux__DOLLAR__515__A),
    .B(__DOLLAR__procmux__DOLLAR__515__B),
    .S(__DOLLAR__procmux__DOLLAR__515__S),
    .Y(__DOLLAR__procmux__DOLLAR__515__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__520' (Module rtMux_U26)
  wire [31:0] __DOLLAR__procmux__DOLLAR__520__A;
  wire [31:0] __DOLLAR__procmux__DOLLAR__520__B;
  wire  __DOLLAR__procmux__DOLLAR__520__S;
  wire [31:0] __DOLLAR__procmux__DOLLAR__520__Y;
  rtMux_U26 __DOLLAR__procmux__DOLLAR__520(
    .A(__DOLLAR__procmux__DOLLAR__520__A),
    .B(__DOLLAR__procmux__DOLLAR__520__B),
    .S(__DOLLAR__procmux__DOLLAR__520__S),
    .Y(__DOLLAR__procmux__DOLLAR__520__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__521_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__521_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__521_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__521_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__521_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__521_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__521_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__522' (Module rtMux_U26)
  wire [31:0] __DOLLAR__procmux__DOLLAR__522__A;
  wire [31:0] __DOLLAR__procmux__DOLLAR__522__B;
  wire  __DOLLAR__procmux__DOLLAR__522__S;
  wire [31:0] __DOLLAR__procmux__DOLLAR__522__Y;
  rtMux_U26 __DOLLAR__procmux__DOLLAR__522(
    .A(__DOLLAR__procmux__DOLLAR__522__A),
    .B(__DOLLAR__procmux__DOLLAR__522__B),
    .S(__DOLLAR__procmux__DOLLAR__522__S),
    .Y(__DOLLAR__procmux__DOLLAR__522__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276(
    .A(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y)
  );

  //All the connections
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__S = __DOLLAR__procmux__DOLLAR__412_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__S = __DOLLAR__procmux__DOLLAR__414_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__S = __DOLLAR__procmux__DOLLAR__417_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__S = __DOLLAR__procmux__DOLLAR__419_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__S = __DOLLAR__procmux__DOLLAR__422_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__S = __DOLLAR__procmux__DOLLAR__424_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__S = __DOLLAR__procmux__DOLLAR__427_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__S = __DOLLAR__procmux__DOLLAR__429_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__S = __DOLLAR__procmux__DOLLAR__432_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__S = __DOLLAR__procmux__DOLLAR__434_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__S = __DOLLAR__procmux__DOLLAR__437_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__S = __DOLLAR__procmux__DOLLAR__439_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__S = __DOLLAR__procmux__DOLLAR__442_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__S = __DOLLAR__procmux__DOLLAR__444_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__S = __DOLLAR__procmux__DOLLAR__447_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__S = __DOLLAR__procmux__DOLLAR__449_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__S = __DOLLAR__procmux__DOLLAR__452_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__S = __DOLLAR__procmux__DOLLAR__454_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__S = __DOLLAR__procmux__DOLLAR__457_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__S = __DOLLAR__procmux__DOLLAR__459_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__S = __DOLLAR__procmux__DOLLAR__462_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__S = __DOLLAR__procmux__DOLLAR__464_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__S = __DOLLAR__procmux__DOLLAR__467_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__S = __DOLLAR__procmux__DOLLAR__469_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__S = __DOLLAR__procmux__DOLLAR__472_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__S = __DOLLAR__procmux__DOLLAR__474_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__S = __DOLLAR__procmux__DOLLAR__477_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__S = __DOLLAR__procmux__DOLLAR__479_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__S = __DOLLAR__procmux__DOLLAR__482_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__S = __DOLLAR__procmux__DOLLAR__484_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__S = __DOLLAR__procmux__DOLLAR__487_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__S = __DOLLAR__procmux__DOLLAR__489_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__S = __DOLLAR__procmux__DOLLAR__492_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__S = __DOLLAR__procmux__DOLLAR__494_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__S = __DOLLAR__procmux__DOLLAR__497_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__S = __DOLLAR__procmux__DOLLAR__499_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__S = __DOLLAR__procmux__DOLLAR__502_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__S = __DOLLAR__procmux__DOLLAR__504_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__S = __DOLLAR__procmux__DOLLAR__507_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__S = __DOLLAR__procmux__DOLLAR__509_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__B[0] = __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procdff__DOLLAR__731__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__731__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__732__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__732__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__733__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__733__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__734__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__734__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__735__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__735__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__736__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__736__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__737__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__737__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__738__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__738__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__739__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__739__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__740__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__740__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__741__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__741__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__742__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__742__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__743__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__743__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__744__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__744__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__745__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__745__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__746__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__746__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__747__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__747__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__748__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__748__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__749__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__749__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__750__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__750__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__751__ARST = reset;
  assign __DOLLAR__procdff__DOLLAR__751__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__412_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__412_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__412_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__413_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__413_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__413_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__414_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__414_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__414_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__415_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__415_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__415_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__417_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__417_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__417_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__418_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__418_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__418_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__419_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__419_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__419_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__420_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__420_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__420_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__422_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__422_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__422_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__423_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__423_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__423_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__424_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__424_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__424_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__425_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__425_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__425_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__427_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__427_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__427_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__428_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__428_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__428_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__429_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__429_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__429_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__430_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__430_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__430_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__432_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__432_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__432_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__433_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__433_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__433_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__434_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__434_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__434_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__435_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__435_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__435_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__437_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__437_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__437_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__438_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__438_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__438_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__439_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__439_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__439_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__440_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__440_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__440_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__442_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__442_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__442_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__443_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__443_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__443_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__444_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__444_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__444_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__445_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__445_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__445_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__447_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__447_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__447_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__448_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__448_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__448_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__449_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__449_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__449_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__450_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__450_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__450_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__452_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__452_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__452_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__453_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__453_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__453_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__454_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__454_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__454_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__455_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__455_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__455_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__457_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__457_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__457_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__458_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__458_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__458_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__459_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__459_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__459_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__460_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__460_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__460_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__462_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__462_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__462_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__463_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__463_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__463_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__464_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__464_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__464_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__465_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__465_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__465_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__467_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__467_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__467_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__468_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__468_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__468_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__469_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__469_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__469_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__470_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__470_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__470_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__472_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__472_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__472_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__473_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__473_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__473_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__474_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__474_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__474_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__475_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__475_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__475_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__477_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__477_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__477_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__478_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__478_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__478_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__479_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__479_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__479_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__480_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__480_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__480_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__482_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__482_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__482_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__483_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__483_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__483_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__484_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__484_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__484_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__485_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__485_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__485_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__487_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__487_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__487_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__488_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__488_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__488_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__489_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__489_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__489_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__490_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__490_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__490_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__492_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__492_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__492_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__493_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__493_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__493_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__494_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__494_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__494_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__495_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__495_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__495_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__497_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__497_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__497_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__498_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__498_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__498_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__499_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__499_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__499_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__500_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__500_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__500_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__502_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__502_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__502_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__503_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__503_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__503_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__504_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__504_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__504_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__505_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__505_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__505_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__507_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__507_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__507_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__508_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__508_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__508_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__509_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__509_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__509_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__510_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__510_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__510_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__513__S = __DOLLAR__procmux__DOLLAR__514_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__514_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__515__S = __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__Y[0];
  assign __DOLLAR__procmux__DOLLAR__520__S = __DOLLAR__procmux__DOLLAR__521_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__521_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__522__S = __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__S = __DOLLAR__procdff__DOLLAR__751__Q[40];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__S = __DOLLAR__procdff__DOLLAR__751__Q[41];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__S = __DOLLAR__procdff__DOLLAR__751__Q[42];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__S = __DOLLAR__procdff__DOLLAR__751__Q[43];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__S = __DOLLAR__procdff__DOLLAR__751__Q[44];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__S = __DOLLAR__procdff__DOLLAR__751__Q[45];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__S = __DOLLAR__procdff__DOLLAR__751__Q[46];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__S = __DOLLAR__procdff__DOLLAR__751__Q[47];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__S = __DOLLAR__procdff__DOLLAR__751__Q[48];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__S = __DOLLAR__procdff__DOLLAR__751__Q[49];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__S = __DOLLAR__procdff__DOLLAR__751__Q[50];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__S = __DOLLAR__procdff__DOLLAR__751__Q[51];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__S = __DOLLAR__procdff__DOLLAR__751__Q[52];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__S = __DOLLAR__procdff__DOLLAR__751__Q[53];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__S = __DOLLAR__procdff__DOLLAR__751__Q[54];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__S = __DOLLAR__procdff__DOLLAR__751__Q[55];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__S = __DOLLAR__procdff__DOLLAR__751__Q[56];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__S = __DOLLAR__procdff__DOLLAR__751__Q[57];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__S = __DOLLAR__procdff__DOLLAR__751__Q[58];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__S = __DOLLAR__procdff__DOLLAR__751__Q[59];
  assign __DOLLAR__eq__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__206__DOLLAR__196__A[0] = config_en;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__A[0] = __DOLLAR__procmux__DOLLAR__413_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__792__B[0] = __DOLLAR__procmux__DOLLAR__412_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__A[0] = __DOLLAR__procmux__DOLLAR__418_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__800__B[0] = __DOLLAR__procmux__DOLLAR__417_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__A[0] = __DOLLAR__procmux__DOLLAR__423_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__808__B[0] = __DOLLAR__procmux__DOLLAR__422_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__A[0] = __DOLLAR__procmux__DOLLAR__428_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__816__B[0] = __DOLLAR__procmux__DOLLAR__427_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__A[0] = __DOLLAR__procmux__DOLLAR__433_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__824__B[0] = __DOLLAR__procmux__DOLLAR__432_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__A[0] = __DOLLAR__procmux__DOLLAR__438_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__832__B[0] = __DOLLAR__procmux__DOLLAR__437_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__A[0] = __DOLLAR__procmux__DOLLAR__443_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__840__B[0] = __DOLLAR__procmux__DOLLAR__442_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__A[0] = __DOLLAR__procmux__DOLLAR__448_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__848__B[0] = __DOLLAR__procmux__DOLLAR__447_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__A[0] = __DOLLAR__procmux__DOLLAR__453_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__856__B[0] = __DOLLAR__procmux__DOLLAR__452_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__A[0] = __DOLLAR__procmux__DOLLAR__458_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__864__B[0] = __DOLLAR__procmux__DOLLAR__457_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__A[0] = __DOLLAR__procmux__DOLLAR__463_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__872__B[0] = __DOLLAR__procmux__DOLLAR__462_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__A[0] = __DOLLAR__procmux__DOLLAR__468_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__880__B[0] = __DOLLAR__procmux__DOLLAR__467_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__A[0] = __DOLLAR__procmux__DOLLAR__473_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__888__B[0] = __DOLLAR__procmux__DOLLAR__472_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__A[0] = __DOLLAR__procmux__DOLLAR__478_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__896__B[0] = __DOLLAR__procmux__DOLLAR__477_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__A[0] = __DOLLAR__procmux__DOLLAR__483_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__904__B[0] = __DOLLAR__procmux__DOLLAR__482_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__A[0] = __DOLLAR__procmux__DOLLAR__488_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__912__B[0] = __DOLLAR__procmux__DOLLAR__487_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__A[0] = __DOLLAR__procmux__DOLLAR__493_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__920__B[0] = __DOLLAR__procmux__DOLLAR__492_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__A[0] = __DOLLAR__procmux__DOLLAR__498_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__928__B[0] = __DOLLAR__procmux__DOLLAR__497_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__A[0] = __DOLLAR__procmux__DOLLAR__503_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__936__B[0] = __DOLLAR__procmux__DOLLAR__502_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__A[0] = __DOLLAR__procmux__DOLLAR__508_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__944__B[0] = __DOLLAR__procmux__DOLLAR__507_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[0] = in_2_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[1] = in_2_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[10] = in_2_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[11] = in_2_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[12] = in_2_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[13] = in_2_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[14] = in_2_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[15] = in_2_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[2] = in_2_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[3] = in_2_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[4] = in_2_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[5] = in_2_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[6] = in_2_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[7] = in_2_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[8] = in_2_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__A[9] = in_2_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__788__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[0] = in_0_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[1] = in_0_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[10] = in_0_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[11] = in_0_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[12] = in_0_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[13] = in_0_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[14] = in_0_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[15] = in_0_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[2] = in_0_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[3] = in_0_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[4] = in_0_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[5] = in_0_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[6] = in_0_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[7] = in_0_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[8] = in_0_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__A[9] = in_0_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[0] = in_1_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[1] = in_1_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[10] = in_1_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[11] = in_1_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[12] = in_1_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[13] = in_1_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[14] = in_1_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[15] = in_1_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[2] = in_1_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[3] = in_1_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[4] = in_1_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[5] = in_1_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[6] = in_1_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[7] = in_1_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[8] = in_1_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__B[9] = in_1_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__790__Y[9];
  assign __DOLLAR__procdff__DOLLAR__731__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[0];
  assign __DOLLAR__procdff__DOLLAR__731__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[1];
  assign __DOLLAR__procdff__DOLLAR__731__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[10];
  assign __DOLLAR__procdff__DOLLAR__731__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[11];
  assign __DOLLAR__procdff__DOLLAR__731__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[12];
  assign __DOLLAR__procdff__DOLLAR__731__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[13];
  assign __DOLLAR__procdff__DOLLAR__731__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[14];
  assign __DOLLAR__procdff__DOLLAR__731__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[15];
  assign __DOLLAR__procdff__DOLLAR__731__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[2];
  assign __DOLLAR__procdff__DOLLAR__731__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[3];
  assign __DOLLAR__procdff__DOLLAR__731__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[4];
  assign __DOLLAR__procdff__DOLLAR__731__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[5];
  assign __DOLLAR__procdff__DOLLAR__731__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[6];
  assign __DOLLAR__procdff__DOLLAR__731__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[7];
  assign __DOLLAR__procdff__DOLLAR__731__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[8];
  assign __DOLLAR__procdff__DOLLAR__731__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__794__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[0] = in_2_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[1] = in_2_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[10] = in_2_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[11] = in_2_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[12] = in_2_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[13] = in_2_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[14] = in_2_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[15] = in_2_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[2] = in_2_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[3] = in_2_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[4] = in_2_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[5] = in_2_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[6] = in_2_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[7] = in_2_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[8] = in_2_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__A[9] = in_2_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__796__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[0] = in_0_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[1] = in_0_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[10] = in_0_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[11] = in_0_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[12] = in_0_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[13] = in_0_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[14] = in_0_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[15] = in_0_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[2] = in_0_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[3] = in_0_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[4] = in_0_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[5] = in_0_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[6] = in_0_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[7] = in_0_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[8] = in_0_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__A[9] = in_0_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[0] = in_1_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[1] = in_1_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[10] = in_1_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[11] = in_1_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[12] = in_1_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[13] = in_1_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[14] = in_1_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[15] = in_1_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[2] = in_1_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[3] = in_1_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[4] = in_1_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[5] = in_1_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[6] = in_1_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[7] = in_1_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[8] = in_1_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__B[9] = in_1_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__798__Y[9];
  assign __DOLLAR__procdff__DOLLAR__732__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[0];
  assign __DOLLAR__procdff__DOLLAR__732__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[1];
  assign __DOLLAR__procdff__DOLLAR__732__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[10];
  assign __DOLLAR__procdff__DOLLAR__732__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[11];
  assign __DOLLAR__procdff__DOLLAR__732__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[12];
  assign __DOLLAR__procdff__DOLLAR__732__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[13];
  assign __DOLLAR__procdff__DOLLAR__732__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[14];
  assign __DOLLAR__procdff__DOLLAR__732__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[15];
  assign __DOLLAR__procdff__DOLLAR__732__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[2];
  assign __DOLLAR__procdff__DOLLAR__732__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[3];
  assign __DOLLAR__procdff__DOLLAR__732__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[4];
  assign __DOLLAR__procdff__DOLLAR__732__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[5];
  assign __DOLLAR__procdff__DOLLAR__732__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[6];
  assign __DOLLAR__procdff__DOLLAR__732__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[7];
  assign __DOLLAR__procdff__DOLLAR__732__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[8];
  assign __DOLLAR__procdff__DOLLAR__732__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__802__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[0] = in_2_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[1] = in_2_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[10] = in_2_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[11] = in_2_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[12] = in_2_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[13] = in_2_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[14] = in_2_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[15] = in_2_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[2] = in_2_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[3] = in_2_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[4] = in_2_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[5] = in_2_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[6] = in_2_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[7] = in_2_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[8] = in_2_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__A[9] = in_2_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__804__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[0] = in_0_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[1] = in_0_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[10] = in_0_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[11] = in_0_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[12] = in_0_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[13] = in_0_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[14] = in_0_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[15] = in_0_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[2] = in_0_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[3] = in_0_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[4] = in_0_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[5] = in_0_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[6] = in_0_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[7] = in_0_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[8] = in_0_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__A[9] = in_0_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[0] = in_1_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[1] = in_1_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[10] = in_1_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[11] = in_1_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[12] = in_1_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[13] = in_1_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[14] = in_1_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[15] = in_1_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[2] = in_1_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[3] = in_1_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[4] = in_1_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[5] = in_1_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[6] = in_1_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[7] = in_1_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[8] = in_1_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__B[9] = in_1_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__806__Y[9];
  assign __DOLLAR__procdff__DOLLAR__733__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[0];
  assign __DOLLAR__procdff__DOLLAR__733__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[1];
  assign __DOLLAR__procdff__DOLLAR__733__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[10];
  assign __DOLLAR__procdff__DOLLAR__733__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[11];
  assign __DOLLAR__procdff__DOLLAR__733__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[12];
  assign __DOLLAR__procdff__DOLLAR__733__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[13];
  assign __DOLLAR__procdff__DOLLAR__733__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[14];
  assign __DOLLAR__procdff__DOLLAR__733__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[15];
  assign __DOLLAR__procdff__DOLLAR__733__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[2];
  assign __DOLLAR__procdff__DOLLAR__733__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[3];
  assign __DOLLAR__procdff__DOLLAR__733__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[4];
  assign __DOLLAR__procdff__DOLLAR__733__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[5];
  assign __DOLLAR__procdff__DOLLAR__733__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[6];
  assign __DOLLAR__procdff__DOLLAR__733__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[7];
  assign __DOLLAR__procdff__DOLLAR__733__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[8];
  assign __DOLLAR__procdff__DOLLAR__733__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__810__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[0] = in_2_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[1] = in_2_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[10] = in_2_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[11] = in_2_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[12] = in_2_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[13] = in_2_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[14] = in_2_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[15] = in_2_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[2] = in_2_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[3] = in_2_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[4] = in_2_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[5] = in_2_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[6] = in_2_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[7] = in_2_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[8] = in_2_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__A[9] = in_2_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__812__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[0] = in_0_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[1] = in_0_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[10] = in_0_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[11] = in_0_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[12] = in_0_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[13] = in_0_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[14] = in_0_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[15] = in_0_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[2] = in_0_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[3] = in_0_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[4] = in_0_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[5] = in_0_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[6] = in_0_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[7] = in_0_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[8] = in_0_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__A[9] = in_0_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[0] = in_1_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[1] = in_1_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[10] = in_1_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[11] = in_1_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[12] = in_1_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[13] = in_1_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[14] = in_1_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[15] = in_1_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[2] = in_1_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[3] = in_1_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[4] = in_1_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[5] = in_1_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[6] = in_1_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[7] = in_1_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[8] = in_1_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__B[9] = in_1_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__814__Y[9];
  assign __DOLLAR__procdff__DOLLAR__734__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[0];
  assign __DOLLAR__procdff__DOLLAR__734__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[1];
  assign __DOLLAR__procdff__DOLLAR__734__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[10];
  assign __DOLLAR__procdff__DOLLAR__734__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[11];
  assign __DOLLAR__procdff__DOLLAR__734__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[12];
  assign __DOLLAR__procdff__DOLLAR__734__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[13];
  assign __DOLLAR__procdff__DOLLAR__734__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[14];
  assign __DOLLAR__procdff__DOLLAR__734__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[15];
  assign __DOLLAR__procdff__DOLLAR__734__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[2];
  assign __DOLLAR__procdff__DOLLAR__734__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[3];
  assign __DOLLAR__procdff__DOLLAR__734__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[4];
  assign __DOLLAR__procdff__DOLLAR__734__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[5];
  assign __DOLLAR__procdff__DOLLAR__734__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[6];
  assign __DOLLAR__procdff__DOLLAR__734__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[7];
  assign __DOLLAR__procdff__DOLLAR__734__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[8];
  assign __DOLLAR__procdff__DOLLAR__734__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__818__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[0] = in_2_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[1] = in_2_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[10] = in_2_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[11] = in_2_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[12] = in_2_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[13] = in_2_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[14] = in_2_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[15] = in_2_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[2] = in_2_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[3] = in_2_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[4] = in_2_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[5] = in_2_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[6] = in_2_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[7] = in_2_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[8] = in_2_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__A[9] = in_2_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__820__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[0] = in_0_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[1] = in_0_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[10] = in_0_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[11] = in_0_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[12] = in_0_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[13] = in_0_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[14] = in_0_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[15] = in_0_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[2] = in_0_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[3] = in_0_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[4] = in_0_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[5] = in_0_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[6] = in_0_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[7] = in_0_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[8] = in_0_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__A[9] = in_0_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[0] = in_1_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[1] = in_1_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[10] = in_1_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[11] = in_1_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[12] = in_1_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[13] = in_1_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[14] = in_1_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[15] = in_1_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[2] = in_1_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[3] = in_1_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[4] = in_1_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[5] = in_1_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[6] = in_1_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[7] = in_1_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[8] = in_1_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__B[9] = in_1_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__822__Y[9];
  assign __DOLLAR__procdff__DOLLAR__735__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[0];
  assign __DOLLAR__procdff__DOLLAR__735__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[1];
  assign __DOLLAR__procdff__DOLLAR__735__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[10];
  assign __DOLLAR__procdff__DOLLAR__735__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[11];
  assign __DOLLAR__procdff__DOLLAR__735__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[12];
  assign __DOLLAR__procdff__DOLLAR__735__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[13];
  assign __DOLLAR__procdff__DOLLAR__735__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[14];
  assign __DOLLAR__procdff__DOLLAR__735__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[15];
  assign __DOLLAR__procdff__DOLLAR__735__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[2];
  assign __DOLLAR__procdff__DOLLAR__735__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[3];
  assign __DOLLAR__procdff__DOLLAR__735__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[4];
  assign __DOLLAR__procdff__DOLLAR__735__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[5];
  assign __DOLLAR__procdff__DOLLAR__735__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[6];
  assign __DOLLAR__procdff__DOLLAR__735__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[7];
  assign __DOLLAR__procdff__DOLLAR__735__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[8];
  assign __DOLLAR__procdff__DOLLAR__735__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__826__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[0] = in_3_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[1] = in_3_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[10] = in_3_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[11] = in_3_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[12] = in_3_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[13] = in_3_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[14] = in_3_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[15] = in_3_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[2] = in_3_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[3] = in_3_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[4] = in_3_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[5] = in_3_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[6] = in_3_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[7] = in_3_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[8] = in_3_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__A[9] = in_3_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__828__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[0] = in_0_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[1] = in_0_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[10] = in_0_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[11] = in_0_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[12] = in_0_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[13] = in_0_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[14] = in_0_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[15] = in_0_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[2] = in_0_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[3] = in_0_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[4] = in_0_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[5] = in_0_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[6] = in_0_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[7] = in_0_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[8] = in_0_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__A[9] = in_0_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[0] = in_1_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[1] = in_1_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[10] = in_1_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[11] = in_1_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[12] = in_1_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[13] = in_1_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[14] = in_1_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[15] = in_1_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[2] = in_1_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[3] = in_1_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[4] = in_1_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[5] = in_1_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[6] = in_1_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[7] = in_1_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[8] = in_1_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__B[9] = in_1_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__830__Y[9];
  assign __DOLLAR__procdff__DOLLAR__736__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[0];
  assign __DOLLAR__procdff__DOLLAR__736__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[1];
  assign __DOLLAR__procdff__DOLLAR__736__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[10];
  assign __DOLLAR__procdff__DOLLAR__736__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[11];
  assign __DOLLAR__procdff__DOLLAR__736__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[12];
  assign __DOLLAR__procdff__DOLLAR__736__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[13];
  assign __DOLLAR__procdff__DOLLAR__736__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[14];
  assign __DOLLAR__procdff__DOLLAR__736__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[15];
  assign __DOLLAR__procdff__DOLLAR__736__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[2];
  assign __DOLLAR__procdff__DOLLAR__736__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[3];
  assign __DOLLAR__procdff__DOLLAR__736__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[4];
  assign __DOLLAR__procdff__DOLLAR__736__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[5];
  assign __DOLLAR__procdff__DOLLAR__736__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[6];
  assign __DOLLAR__procdff__DOLLAR__736__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[7];
  assign __DOLLAR__procdff__DOLLAR__736__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[8];
  assign __DOLLAR__procdff__DOLLAR__736__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__834__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[0] = in_3_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[1] = in_3_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[10] = in_3_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[11] = in_3_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[12] = in_3_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[13] = in_3_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[14] = in_3_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[15] = in_3_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[2] = in_3_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[3] = in_3_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[4] = in_3_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[5] = in_3_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[6] = in_3_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[7] = in_3_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[8] = in_3_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__A[9] = in_3_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__836__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[0] = in_0_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[1] = in_0_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[10] = in_0_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[11] = in_0_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[12] = in_0_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[13] = in_0_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[14] = in_0_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[15] = in_0_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[2] = in_0_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[3] = in_0_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[4] = in_0_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[5] = in_0_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[6] = in_0_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[7] = in_0_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[8] = in_0_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__A[9] = in_0_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[0] = in_1_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[1] = in_1_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[10] = in_1_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[11] = in_1_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[12] = in_1_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[13] = in_1_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[14] = in_1_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[15] = in_1_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[2] = in_1_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[3] = in_1_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[4] = in_1_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[5] = in_1_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[6] = in_1_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[7] = in_1_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[8] = in_1_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__B[9] = in_1_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__838__Y[9];
  assign __DOLLAR__procdff__DOLLAR__737__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[0];
  assign __DOLLAR__procdff__DOLLAR__737__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[1];
  assign __DOLLAR__procdff__DOLLAR__737__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[10];
  assign __DOLLAR__procdff__DOLLAR__737__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[11];
  assign __DOLLAR__procdff__DOLLAR__737__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[12];
  assign __DOLLAR__procdff__DOLLAR__737__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[13];
  assign __DOLLAR__procdff__DOLLAR__737__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[14];
  assign __DOLLAR__procdff__DOLLAR__737__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[15];
  assign __DOLLAR__procdff__DOLLAR__737__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[2];
  assign __DOLLAR__procdff__DOLLAR__737__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[3];
  assign __DOLLAR__procdff__DOLLAR__737__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[4];
  assign __DOLLAR__procdff__DOLLAR__737__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[5];
  assign __DOLLAR__procdff__DOLLAR__737__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[6];
  assign __DOLLAR__procdff__DOLLAR__737__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[7];
  assign __DOLLAR__procdff__DOLLAR__737__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[8];
  assign __DOLLAR__procdff__DOLLAR__737__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__842__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[0] = in_3_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[1] = in_3_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[10] = in_3_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[11] = in_3_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[12] = in_3_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[13] = in_3_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[14] = in_3_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[15] = in_3_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[2] = in_3_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[3] = in_3_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[4] = in_3_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[5] = in_3_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[6] = in_3_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[7] = in_3_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[8] = in_3_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__A[9] = in_3_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__844__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[0] = in_0_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[1] = in_0_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[10] = in_0_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[11] = in_0_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[12] = in_0_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[13] = in_0_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[14] = in_0_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[15] = in_0_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[2] = in_0_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[3] = in_0_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[4] = in_0_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[5] = in_0_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[6] = in_0_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[7] = in_0_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[8] = in_0_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__A[9] = in_0_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[0] = in_1_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[1] = in_1_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[10] = in_1_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[11] = in_1_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[12] = in_1_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[13] = in_1_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[14] = in_1_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[15] = in_1_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[2] = in_1_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[3] = in_1_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[4] = in_1_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[5] = in_1_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[6] = in_1_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[7] = in_1_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[8] = in_1_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__B[9] = in_1_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__846__Y[9];
  assign __DOLLAR__procdff__DOLLAR__738__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[0];
  assign __DOLLAR__procdff__DOLLAR__738__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[1];
  assign __DOLLAR__procdff__DOLLAR__738__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[10];
  assign __DOLLAR__procdff__DOLLAR__738__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[11];
  assign __DOLLAR__procdff__DOLLAR__738__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[12];
  assign __DOLLAR__procdff__DOLLAR__738__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[13];
  assign __DOLLAR__procdff__DOLLAR__738__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[14];
  assign __DOLLAR__procdff__DOLLAR__738__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[15];
  assign __DOLLAR__procdff__DOLLAR__738__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[2];
  assign __DOLLAR__procdff__DOLLAR__738__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[3];
  assign __DOLLAR__procdff__DOLLAR__738__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[4];
  assign __DOLLAR__procdff__DOLLAR__738__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[5];
  assign __DOLLAR__procdff__DOLLAR__738__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[6];
  assign __DOLLAR__procdff__DOLLAR__738__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[7];
  assign __DOLLAR__procdff__DOLLAR__738__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[8];
  assign __DOLLAR__procdff__DOLLAR__738__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__850__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[0] = in_3_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[1] = in_3_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[10] = in_3_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[11] = in_3_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[12] = in_3_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[13] = in_3_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[14] = in_3_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[15] = in_3_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[2] = in_3_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[3] = in_3_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[4] = in_3_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[5] = in_3_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[6] = in_3_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[7] = in_3_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[8] = in_3_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__A[9] = in_3_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__852__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[0] = in_0_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[1] = in_0_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[10] = in_0_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[11] = in_0_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[12] = in_0_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[13] = in_0_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[14] = in_0_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[15] = in_0_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[2] = in_0_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[3] = in_0_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[4] = in_0_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[5] = in_0_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[6] = in_0_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[7] = in_0_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[8] = in_0_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__A[9] = in_0_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[0] = in_1_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[1] = in_1_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[10] = in_1_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[11] = in_1_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[12] = in_1_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[13] = in_1_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[14] = in_1_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[15] = in_1_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[2] = in_1_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[3] = in_1_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[4] = in_1_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[5] = in_1_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[6] = in_1_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[7] = in_1_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[8] = in_1_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__B[9] = in_1_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__854__Y[9];
  assign __DOLLAR__procdff__DOLLAR__739__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[0];
  assign __DOLLAR__procdff__DOLLAR__739__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[1];
  assign __DOLLAR__procdff__DOLLAR__739__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[10];
  assign __DOLLAR__procdff__DOLLAR__739__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[11];
  assign __DOLLAR__procdff__DOLLAR__739__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[12];
  assign __DOLLAR__procdff__DOLLAR__739__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[13];
  assign __DOLLAR__procdff__DOLLAR__739__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[14];
  assign __DOLLAR__procdff__DOLLAR__739__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[15];
  assign __DOLLAR__procdff__DOLLAR__739__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[2];
  assign __DOLLAR__procdff__DOLLAR__739__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[3];
  assign __DOLLAR__procdff__DOLLAR__739__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[4];
  assign __DOLLAR__procdff__DOLLAR__739__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[5];
  assign __DOLLAR__procdff__DOLLAR__739__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[6];
  assign __DOLLAR__procdff__DOLLAR__739__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[7];
  assign __DOLLAR__procdff__DOLLAR__739__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[8];
  assign __DOLLAR__procdff__DOLLAR__739__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__858__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[0] = in_3_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[1] = in_3_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[10] = in_3_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[11] = in_3_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[12] = in_3_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[13] = in_3_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[14] = in_3_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[15] = in_3_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[2] = in_3_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[3] = in_3_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[4] = in_3_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[5] = in_3_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[6] = in_3_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[7] = in_3_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[8] = in_3_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__A[9] = in_3_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__860__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[0] = in_0_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[1] = in_0_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[10] = in_0_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[11] = in_0_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[12] = in_0_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[13] = in_0_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[14] = in_0_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[15] = in_0_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[2] = in_0_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[3] = in_0_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[4] = in_0_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[5] = in_0_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[6] = in_0_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[7] = in_0_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[8] = in_0_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__A[9] = in_0_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[0] = in_1_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[1] = in_1_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[10] = in_1_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[11] = in_1_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[12] = in_1_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[13] = in_1_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[14] = in_1_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[15] = in_1_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[2] = in_1_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[3] = in_1_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[4] = in_1_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[5] = in_1_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[6] = in_1_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[7] = in_1_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[8] = in_1_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__B[9] = in_1_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__862__Y[9];
  assign __DOLLAR__procdff__DOLLAR__740__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[0];
  assign __DOLLAR__procdff__DOLLAR__740__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[1];
  assign __DOLLAR__procdff__DOLLAR__740__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[10];
  assign __DOLLAR__procdff__DOLLAR__740__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[11];
  assign __DOLLAR__procdff__DOLLAR__740__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[12];
  assign __DOLLAR__procdff__DOLLAR__740__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[13];
  assign __DOLLAR__procdff__DOLLAR__740__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[14];
  assign __DOLLAR__procdff__DOLLAR__740__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[15];
  assign __DOLLAR__procdff__DOLLAR__740__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[2];
  assign __DOLLAR__procdff__DOLLAR__740__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[3];
  assign __DOLLAR__procdff__DOLLAR__740__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[4];
  assign __DOLLAR__procdff__DOLLAR__740__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[5];
  assign __DOLLAR__procdff__DOLLAR__740__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[6];
  assign __DOLLAR__procdff__DOLLAR__740__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[7];
  assign __DOLLAR__procdff__DOLLAR__740__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[8];
  assign __DOLLAR__procdff__DOLLAR__740__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__866__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[0] = in_3_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[1] = in_3_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[10] = in_3_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[11] = in_3_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[12] = in_3_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[13] = in_3_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[14] = in_3_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[15] = in_3_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[2] = in_3_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[3] = in_3_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[4] = in_3_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[5] = in_3_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[6] = in_3_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[7] = in_3_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[8] = in_3_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__A[9] = in_3_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__868__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[0] = in_0_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[1] = in_0_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[10] = in_0_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[11] = in_0_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[12] = in_0_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[13] = in_0_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[14] = in_0_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[15] = in_0_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[2] = in_0_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[3] = in_0_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[4] = in_0_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[5] = in_0_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[6] = in_0_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[7] = in_0_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[8] = in_0_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__A[9] = in_0_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[0] = in_2_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[1] = in_2_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[10] = in_2_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[11] = in_2_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[12] = in_2_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[13] = in_2_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[14] = in_2_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[15] = in_2_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[2] = in_2_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[3] = in_2_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[4] = in_2_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[5] = in_2_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[6] = in_2_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[7] = in_2_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[8] = in_2_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__B[9] = in_2_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__870__Y[9];
  assign __DOLLAR__procdff__DOLLAR__741__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[0];
  assign __DOLLAR__procdff__DOLLAR__741__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[1];
  assign __DOLLAR__procdff__DOLLAR__741__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[10];
  assign __DOLLAR__procdff__DOLLAR__741__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[11];
  assign __DOLLAR__procdff__DOLLAR__741__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[12];
  assign __DOLLAR__procdff__DOLLAR__741__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[13];
  assign __DOLLAR__procdff__DOLLAR__741__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[14];
  assign __DOLLAR__procdff__DOLLAR__741__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[15];
  assign __DOLLAR__procdff__DOLLAR__741__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[2];
  assign __DOLLAR__procdff__DOLLAR__741__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[3];
  assign __DOLLAR__procdff__DOLLAR__741__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[4];
  assign __DOLLAR__procdff__DOLLAR__741__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[5];
  assign __DOLLAR__procdff__DOLLAR__741__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[6];
  assign __DOLLAR__procdff__DOLLAR__741__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[7];
  assign __DOLLAR__procdff__DOLLAR__741__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[8];
  assign __DOLLAR__procdff__DOLLAR__741__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__874__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[0] = in_3_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[1] = in_3_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[10] = in_3_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[11] = in_3_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[12] = in_3_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[13] = in_3_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[14] = in_3_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[15] = in_3_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[2] = in_3_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[3] = in_3_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[4] = in_3_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[5] = in_3_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[6] = in_3_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[7] = in_3_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[8] = in_3_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__A[9] = in_3_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__876__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[0] = in_0_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[1] = in_0_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[10] = in_0_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[11] = in_0_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[12] = in_0_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[13] = in_0_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[14] = in_0_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[15] = in_0_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[2] = in_0_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[3] = in_0_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[4] = in_0_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[5] = in_0_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[6] = in_0_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[7] = in_0_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[8] = in_0_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__A[9] = in_0_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[0] = in_2_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[1] = in_2_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[10] = in_2_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[11] = in_2_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[12] = in_2_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[13] = in_2_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[14] = in_2_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[15] = in_2_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[2] = in_2_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[3] = in_2_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[4] = in_2_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[5] = in_2_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[6] = in_2_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[7] = in_2_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[8] = in_2_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__B[9] = in_2_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__878__Y[9];
  assign __DOLLAR__procdff__DOLLAR__742__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[0];
  assign __DOLLAR__procdff__DOLLAR__742__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[1];
  assign __DOLLAR__procdff__DOLLAR__742__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[10];
  assign __DOLLAR__procdff__DOLLAR__742__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[11];
  assign __DOLLAR__procdff__DOLLAR__742__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[12];
  assign __DOLLAR__procdff__DOLLAR__742__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[13];
  assign __DOLLAR__procdff__DOLLAR__742__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[14];
  assign __DOLLAR__procdff__DOLLAR__742__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[15];
  assign __DOLLAR__procdff__DOLLAR__742__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[2];
  assign __DOLLAR__procdff__DOLLAR__742__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[3];
  assign __DOLLAR__procdff__DOLLAR__742__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[4];
  assign __DOLLAR__procdff__DOLLAR__742__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[5];
  assign __DOLLAR__procdff__DOLLAR__742__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[6];
  assign __DOLLAR__procdff__DOLLAR__742__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[7];
  assign __DOLLAR__procdff__DOLLAR__742__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[8];
  assign __DOLLAR__procdff__DOLLAR__742__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__882__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[0] = in_3_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[1] = in_3_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[10] = in_3_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[11] = in_3_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[12] = in_3_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[13] = in_3_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[14] = in_3_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[15] = in_3_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[2] = in_3_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[3] = in_3_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[4] = in_3_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[5] = in_3_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[6] = in_3_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[7] = in_3_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[8] = in_3_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__A[9] = in_3_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__884__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[0] = in_0_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[1] = in_0_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[10] = in_0_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[11] = in_0_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[12] = in_0_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[13] = in_0_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[14] = in_0_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[15] = in_0_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[2] = in_0_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[3] = in_0_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[4] = in_0_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[5] = in_0_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[6] = in_0_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[7] = in_0_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[8] = in_0_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__A[9] = in_0_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[0] = in_2_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[1] = in_2_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[10] = in_2_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[11] = in_2_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[12] = in_2_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[13] = in_2_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[14] = in_2_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[15] = in_2_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[2] = in_2_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[3] = in_2_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[4] = in_2_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[5] = in_2_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[6] = in_2_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[7] = in_2_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[8] = in_2_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__B[9] = in_2_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__886__Y[9];
  assign __DOLLAR__procdff__DOLLAR__743__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[0];
  assign __DOLLAR__procdff__DOLLAR__743__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[1];
  assign __DOLLAR__procdff__DOLLAR__743__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[10];
  assign __DOLLAR__procdff__DOLLAR__743__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[11];
  assign __DOLLAR__procdff__DOLLAR__743__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[12];
  assign __DOLLAR__procdff__DOLLAR__743__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[13];
  assign __DOLLAR__procdff__DOLLAR__743__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[14];
  assign __DOLLAR__procdff__DOLLAR__743__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[15];
  assign __DOLLAR__procdff__DOLLAR__743__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[2];
  assign __DOLLAR__procdff__DOLLAR__743__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[3];
  assign __DOLLAR__procdff__DOLLAR__743__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[4];
  assign __DOLLAR__procdff__DOLLAR__743__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[5];
  assign __DOLLAR__procdff__DOLLAR__743__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[6];
  assign __DOLLAR__procdff__DOLLAR__743__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[7];
  assign __DOLLAR__procdff__DOLLAR__743__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[8];
  assign __DOLLAR__procdff__DOLLAR__743__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__890__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[0] = in_3_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[1] = in_3_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[10] = in_3_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[11] = in_3_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[12] = in_3_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[13] = in_3_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[14] = in_3_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[15] = in_3_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[2] = in_3_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[3] = in_3_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[4] = in_3_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[5] = in_3_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[6] = in_3_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[7] = in_3_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[8] = in_3_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__A[9] = in_3_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__892__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[0] = in_0_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[1] = in_0_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[10] = in_0_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[11] = in_0_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[12] = in_0_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[13] = in_0_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[14] = in_0_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[15] = in_0_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[2] = in_0_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[3] = in_0_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[4] = in_0_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[5] = in_0_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[6] = in_0_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[7] = in_0_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[8] = in_0_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__A[9] = in_0_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[0] = in_2_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[1] = in_2_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[10] = in_2_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[11] = in_2_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[12] = in_2_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[13] = in_2_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[14] = in_2_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[15] = in_2_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[2] = in_2_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[3] = in_2_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[4] = in_2_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[5] = in_2_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[6] = in_2_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[7] = in_2_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[8] = in_2_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__B[9] = in_2_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__894__Y[9];
  assign __DOLLAR__procdff__DOLLAR__744__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[0];
  assign __DOLLAR__procdff__DOLLAR__744__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[1];
  assign __DOLLAR__procdff__DOLLAR__744__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[10];
  assign __DOLLAR__procdff__DOLLAR__744__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[11];
  assign __DOLLAR__procdff__DOLLAR__744__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[12];
  assign __DOLLAR__procdff__DOLLAR__744__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[13];
  assign __DOLLAR__procdff__DOLLAR__744__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[14];
  assign __DOLLAR__procdff__DOLLAR__744__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[15];
  assign __DOLLAR__procdff__DOLLAR__744__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[2];
  assign __DOLLAR__procdff__DOLLAR__744__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[3];
  assign __DOLLAR__procdff__DOLLAR__744__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[4];
  assign __DOLLAR__procdff__DOLLAR__744__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[5];
  assign __DOLLAR__procdff__DOLLAR__744__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[6];
  assign __DOLLAR__procdff__DOLLAR__744__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[7];
  assign __DOLLAR__procdff__DOLLAR__744__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[8];
  assign __DOLLAR__procdff__DOLLAR__744__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__898__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[0] = in_3_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[1] = in_3_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[10] = in_3_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[11] = in_3_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[12] = in_3_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[13] = in_3_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[14] = in_3_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[15] = in_3_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[2] = in_3_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[3] = in_3_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[4] = in_3_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[5] = in_3_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[6] = in_3_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[7] = in_3_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[8] = in_3_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__A[9] = in_3_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__900__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[0] = in_0_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[1] = in_0_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[10] = in_0_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[11] = in_0_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[12] = in_0_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[13] = in_0_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[14] = in_0_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[15] = in_0_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[2] = in_0_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[3] = in_0_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[4] = in_0_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[5] = in_0_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[6] = in_0_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[7] = in_0_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[8] = in_0_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__A[9] = in_0_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[0] = in_2_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[1] = in_2_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[10] = in_2_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[11] = in_2_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[12] = in_2_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[13] = in_2_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[14] = in_2_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[15] = in_2_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[2] = in_2_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[3] = in_2_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[4] = in_2_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[5] = in_2_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[6] = in_2_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[7] = in_2_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[8] = in_2_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__B[9] = in_2_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__902__Y[9];
  assign __DOLLAR__procdff__DOLLAR__745__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[0];
  assign __DOLLAR__procdff__DOLLAR__745__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[1];
  assign __DOLLAR__procdff__DOLLAR__745__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[10];
  assign __DOLLAR__procdff__DOLLAR__745__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[11];
  assign __DOLLAR__procdff__DOLLAR__745__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[12];
  assign __DOLLAR__procdff__DOLLAR__745__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[13];
  assign __DOLLAR__procdff__DOLLAR__745__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[14];
  assign __DOLLAR__procdff__DOLLAR__745__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[15];
  assign __DOLLAR__procdff__DOLLAR__745__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[2];
  assign __DOLLAR__procdff__DOLLAR__745__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[3];
  assign __DOLLAR__procdff__DOLLAR__745__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[4];
  assign __DOLLAR__procdff__DOLLAR__745__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[5];
  assign __DOLLAR__procdff__DOLLAR__745__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[6];
  assign __DOLLAR__procdff__DOLLAR__745__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[7];
  assign __DOLLAR__procdff__DOLLAR__745__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[8];
  assign __DOLLAR__procdff__DOLLAR__745__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__906__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[0] = in_3_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[1] = in_3_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[10] = in_3_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[11] = in_3_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[12] = in_3_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[13] = in_3_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[14] = in_3_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[15] = in_3_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[2] = in_3_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[3] = in_3_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[4] = in_3_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[5] = in_3_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[6] = in_3_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[7] = in_3_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[8] = in_3_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__A[9] = in_3_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__908__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[0] = in_1_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[1] = in_1_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[10] = in_1_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[11] = in_1_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[12] = in_1_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[13] = in_1_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[14] = in_1_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[15] = in_1_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[2] = in_1_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[3] = in_1_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[4] = in_1_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[5] = in_1_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[6] = in_1_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[7] = in_1_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[8] = in_1_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__A[9] = in_1_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[0] = in_2_4[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[1] = in_2_4[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[10] = in_2_4[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[11] = in_2_4[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[12] = in_2_4[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[13] = in_2_4[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[14] = in_2_4[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[15] = in_2_4[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[2] = in_2_4[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[3] = in_2_4[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[4] = in_2_4[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[5] = in_2_4[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[6] = in_2_4[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[7] = in_2_4[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[8] = in_2_4[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__B[9] = in_2_4[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__910__Y[9];
  assign __DOLLAR__procdff__DOLLAR__746__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[0];
  assign __DOLLAR__procdff__DOLLAR__746__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[1];
  assign __DOLLAR__procdff__DOLLAR__746__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[10];
  assign __DOLLAR__procdff__DOLLAR__746__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[11];
  assign __DOLLAR__procdff__DOLLAR__746__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[12];
  assign __DOLLAR__procdff__DOLLAR__746__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[13];
  assign __DOLLAR__procdff__DOLLAR__746__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[14];
  assign __DOLLAR__procdff__DOLLAR__746__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[15];
  assign __DOLLAR__procdff__DOLLAR__746__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[2];
  assign __DOLLAR__procdff__DOLLAR__746__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[3];
  assign __DOLLAR__procdff__DOLLAR__746__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[4];
  assign __DOLLAR__procdff__DOLLAR__746__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[5];
  assign __DOLLAR__procdff__DOLLAR__746__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[6];
  assign __DOLLAR__procdff__DOLLAR__746__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[7];
  assign __DOLLAR__procdff__DOLLAR__746__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[8];
  assign __DOLLAR__procdff__DOLLAR__746__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__914__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[0] = in_3_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[1] = in_3_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[10] = in_3_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[11] = in_3_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[12] = in_3_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[13] = in_3_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[14] = in_3_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[15] = in_3_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[2] = in_3_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[3] = in_3_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[4] = in_3_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[5] = in_3_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[6] = in_3_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[7] = in_3_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[8] = in_3_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__A[9] = in_3_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__916__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[0] = in_1_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[1] = in_1_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[10] = in_1_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[11] = in_1_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[12] = in_1_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[13] = in_1_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[14] = in_1_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[15] = in_1_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[2] = in_1_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[3] = in_1_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[4] = in_1_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[5] = in_1_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[6] = in_1_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[7] = in_1_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[8] = in_1_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__A[9] = in_1_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[0] = in_2_3[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[1] = in_2_3[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[10] = in_2_3[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[11] = in_2_3[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[12] = in_2_3[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[13] = in_2_3[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[14] = in_2_3[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[15] = in_2_3[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[2] = in_2_3[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[3] = in_2_3[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[4] = in_2_3[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[5] = in_2_3[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[6] = in_2_3[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[7] = in_2_3[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[8] = in_2_3[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__B[9] = in_2_3[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__918__Y[9];
  assign __DOLLAR__procdff__DOLLAR__747__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[0];
  assign __DOLLAR__procdff__DOLLAR__747__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[1];
  assign __DOLLAR__procdff__DOLLAR__747__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[10];
  assign __DOLLAR__procdff__DOLLAR__747__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[11];
  assign __DOLLAR__procdff__DOLLAR__747__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[12];
  assign __DOLLAR__procdff__DOLLAR__747__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[13];
  assign __DOLLAR__procdff__DOLLAR__747__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[14];
  assign __DOLLAR__procdff__DOLLAR__747__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[15];
  assign __DOLLAR__procdff__DOLLAR__747__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[2];
  assign __DOLLAR__procdff__DOLLAR__747__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[3];
  assign __DOLLAR__procdff__DOLLAR__747__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[4];
  assign __DOLLAR__procdff__DOLLAR__747__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[5];
  assign __DOLLAR__procdff__DOLLAR__747__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[6];
  assign __DOLLAR__procdff__DOLLAR__747__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[7];
  assign __DOLLAR__procdff__DOLLAR__747__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[8];
  assign __DOLLAR__procdff__DOLLAR__747__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__922__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[0] = in_3_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[1] = in_3_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[10] = in_3_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[11] = in_3_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[12] = in_3_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[13] = in_3_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[14] = in_3_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[15] = in_3_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[2] = in_3_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[3] = in_3_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[4] = in_3_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[5] = in_3_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[6] = in_3_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[7] = in_3_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[8] = in_3_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__A[9] = in_3_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__924__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[0] = in_1_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[1] = in_1_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[10] = in_1_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[11] = in_1_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[12] = in_1_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[13] = in_1_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[14] = in_1_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[15] = in_1_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[2] = in_1_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[3] = in_1_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[4] = in_1_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[5] = in_1_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[6] = in_1_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[7] = in_1_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[8] = in_1_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__A[9] = in_1_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[0] = in_2_2[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[1] = in_2_2[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[10] = in_2_2[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[11] = in_2_2[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[12] = in_2_2[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[13] = in_2_2[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[14] = in_2_2[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[15] = in_2_2[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[2] = in_2_2[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[3] = in_2_2[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[4] = in_2_2[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[5] = in_2_2[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[6] = in_2_2[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[7] = in_2_2[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[8] = in_2_2[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__B[9] = in_2_2[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__926__Y[9];
  assign __DOLLAR__procdff__DOLLAR__748__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[0];
  assign __DOLLAR__procdff__DOLLAR__748__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[1];
  assign __DOLLAR__procdff__DOLLAR__748__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[10];
  assign __DOLLAR__procdff__DOLLAR__748__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[11];
  assign __DOLLAR__procdff__DOLLAR__748__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[12];
  assign __DOLLAR__procdff__DOLLAR__748__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[13];
  assign __DOLLAR__procdff__DOLLAR__748__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[14];
  assign __DOLLAR__procdff__DOLLAR__748__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[15];
  assign __DOLLAR__procdff__DOLLAR__748__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[2];
  assign __DOLLAR__procdff__DOLLAR__748__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[3];
  assign __DOLLAR__procdff__DOLLAR__748__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[4];
  assign __DOLLAR__procdff__DOLLAR__748__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[5];
  assign __DOLLAR__procdff__DOLLAR__748__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[6];
  assign __DOLLAR__procdff__DOLLAR__748__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[7];
  assign __DOLLAR__procdff__DOLLAR__748__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[8];
  assign __DOLLAR__procdff__DOLLAR__748__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__930__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[0] = in_3_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[1] = in_3_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[10] = in_3_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[11] = in_3_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[12] = in_3_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[13] = in_3_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[14] = in_3_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[15] = in_3_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[2] = in_3_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[3] = in_3_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[4] = in_3_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[5] = in_3_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[6] = in_3_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[7] = in_3_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[8] = in_3_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__A[9] = in_3_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__932__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[0] = in_1_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[1] = in_1_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[10] = in_1_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[11] = in_1_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[12] = in_1_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[13] = in_1_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[14] = in_1_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[15] = in_1_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[2] = in_1_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[3] = in_1_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[4] = in_1_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[5] = in_1_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[6] = in_1_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[7] = in_1_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[8] = in_1_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__A[9] = in_1_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[0] = in_2_1[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[1] = in_2_1[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[10] = in_2_1[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[11] = in_2_1[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[12] = in_2_1[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[13] = in_2_1[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[14] = in_2_1[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[15] = in_2_1[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[2] = in_2_1[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[3] = in_2_1[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[4] = in_2_1[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[5] = in_2_1[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[6] = in_2_1[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[7] = in_2_1[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[8] = in_2_1[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__B[9] = in_2_1[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__934__Y[9];
  assign __DOLLAR__procdff__DOLLAR__749__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[0];
  assign __DOLLAR__procdff__DOLLAR__749__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[1];
  assign __DOLLAR__procdff__DOLLAR__749__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[10];
  assign __DOLLAR__procdff__DOLLAR__749__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[11];
  assign __DOLLAR__procdff__DOLLAR__749__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[12];
  assign __DOLLAR__procdff__DOLLAR__749__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[13];
  assign __DOLLAR__procdff__DOLLAR__749__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[14];
  assign __DOLLAR__procdff__DOLLAR__749__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[15];
  assign __DOLLAR__procdff__DOLLAR__749__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[2];
  assign __DOLLAR__procdff__DOLLAR__749__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[3];
  assign __DOLLAR__procdff__DOLLAR__749__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[4];
  assign __DOLLAR__procdff__DOLLAR__749__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[5];
  assign __DOLLAR__procdff__DOLLAR__749__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[6];
  assign __DOLLAR__procdff__DOLLAR__749__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[7];
  assign __DOLLAR__procdff__DOLLAR__749__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[8];
  assign __DOLLAR__procdff__DOLLAR__749__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__938__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[0] = in_3_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[1] = in_3_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[10] = in_3_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[11] = in_3_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[12] = in_3_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[13] = in_3_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[14] = in_3_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[15] = in_3_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[2] = in_3_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[3] = in_3_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[4] = in_3_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[5] = in_3_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[6] = in_3_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[7] = in_3_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[8] = in_3_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__A[9] = in_3_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[0] = pe_output_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[1] = pe_output_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[10] = pe_output_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[11] = pe_output_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[12] = pe_output_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[13] = pe_output_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[14] = pe_output_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[15] = pe_output_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[2] = pe_output_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[3] = pe_output_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[4] = pe_output_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[5] = pe_output_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[6] = pe_output_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[7] = pe_output_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[8] = pe_output_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__B[9] = pe_output_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__940__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[0] = in_1_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[1] = in_1_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[10] = in_1_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[11] = in_1_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[12] = in_1_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[13] = in_1_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[14] = in_1_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[15] = in_1_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[2] = in_1_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[3] = in_1_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[4] = in_1_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[5] = in_1_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[6] = in_1_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[7] = in_1_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[8] = in_1_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__A[9] = in_1_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[0] = in_2_0[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[1] = in_2_0[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[10] = in_2_0[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[11] = in_2_0[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[12] = in_2_0[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[13] = in_2_0[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[14] = in_2_0[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[15] = in_2_0[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[2] = in_2_0[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[3] = in_2_0[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[4] = in_2_0[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[5] = in_2_0[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[6] = in_2_0[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[7] = in_2_0[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[8] = in_2_0[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__B[9] = in_2_0[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__942__Y[9];
  assign __DOLLAR__procdff__DOLLAR__750__D[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[0];
  assign __DOLLAR__procdff__DOLLAR__750__D[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[1];
  assign __DOLLAR__procdff__DOLLAR__750__D[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[10];
  assign __DOLLAR__procdff__DOLLAR__750__D[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[11];
  assign __DOLLAR__procdff__DOLLAR__750__D[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[12];
  assign __DOLLAR__procdff__DOLLAR__750__D[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[13];
  assign __DOLLAR__procdff__DOLLAR__750__D[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[14];
  assign __DOLLAR__procdff__DOLLAR__750__D[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[15];
  assign __DOLLAR__procdff__DOLLAR__750__D[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[2];
  assign __DOLLAR__procdff__DOLLAR__750__D[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[3];
  assign __DOLLAR__procdff__DOLLAR__750__D[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[4];
  assign __DOLLAR__procdff__DOLLAR__750__D[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[5];
  assign __DOLLAR__procdff__DOLLAR__750__D[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[6];
  assign __DOLLAR__procdff__DOLLAR__750__D[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[7];
  assign __DOLLAR__procdff__DOLLAR__750__D[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[8];
  assign __DOLLAR__procdff__DOLLAR__750__D[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__946__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[0] = __DOLLAR__procdff__DOLLAR__731__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[1] = __DOLLAR__procdff__DOLLAR__731__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[10] = __DOLLAR__procdff__DOLLAR__731__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[11] = __DOLLAR__procdff__DOLLAR__731__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[12] = __DOLLAR__procdff__DOLLAR__731__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[13] = __DOLLAR__procdff__DOLLAR__731__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[14] = __DOLLAR__procdff__DOLLAR__731__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[15] = __DOLLAR__procdff__DOLLAR__731__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[2] = __DOLLAR__procdff__DOLLAR__731__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[3] = __DOLLAR__procdff__DOLLAR__731__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[4] = __DOLLAR__procdff__DOLLAR__731__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[5] = __DOLLAR__procdff__DOLLAR__731__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[6] = __DOLLAR__procdff__DOLLAR__731__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[7] = __DOLLAR__procdff__DOLLAR__731__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[8] = __DOLLAR__procdff__DOLLAR__731__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__B[9] = __DOLLAR__procdff__DOLLAR__731__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[0] = __DOLLAR__procdff__DOLLAR__732__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[1] = __DOLLAR__procdff__DOLLAR__732__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[10] = __DOLLAR__procdff__DOLLAR__732__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[11] = __DOLLAR__procdff__DOLLAR__732__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[12] = __DOLLAR__procdff__DOLLAR__732__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[13] = __DOLLAR__procdff__DOLLAR__732__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[14] = __DOLLAR__procdff__DOLLAR__732__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[15] = __DOLLAR__procdff__DOLLAR__732__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[2] = __DOLLAR__procdff__DOLLAR__732__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[3] = __DOLLAR__procdff__DOLLAR__732__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[4] = __DOLLAR__procdff__DOLLAR__732__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[5] = __DOLLAR__procdff__DOLLAR__732__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[6] = __DOLLAR__procdff__DOLLAR__732__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[7] = __DOLLAR__procdff__DOLLAR__732__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[8] = __DOLLAR__procdff__DOLLAR__732__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__B[9] = __DOLLAR__procdff__DOLLAR__732__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[0] = __DOLLAR__procdff__DOLLAR__733__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[1] = __DOLLAR__procdff__DOLLAR__733__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[10] = __DOLLAR__procdff__DOLLAR__733__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[11] = __DOLLAR__procdff__DOLLAR__733__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[12] = __DOLLAR__procdff__DOLLAR__733__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[13] = __DOLLAR__procdff__DOLLAR__733__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[14] = __DOLLAR__procdff__DOLLAR__733__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[15] = __DOLLAR__procdff__DOLLAR__733__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[2] = __DOLLAR__procdff__DOLLAR__733__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[3] = __DOLLAR__procdff__DOLLAR__733__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[4] = __DOLLAR__procdff__DOLLAR__733__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[5] = __DOLLAR__procdff__DOLLAR__733__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[6] = __DOLLAR__procdff__DOLLAR__733__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[7] = __DOLLAR__procdff__DOLLAR__733__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[8] = __DOLLAR__procdff__DOLLAR__733__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__B[9] = __DOLLAR__procdff__DOLLAR__733__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[0] = __DOLLAR__procdff__DOLLAR__734__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[1] = __DOLLAR__procdff__DOLLAR__734__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[10] = __DOLLAR__procdff__DOLLAR__734__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[11] = __DOLLAR__procdff__DOLLAR__734__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[12] = __DOLLAR__procdff__DOLLAR__734__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[13] = __DOLLAR__procdff__DOLLAR__734__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[14] = __DOLLAR__procdff__DOLLAR__734__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[15] = __DOLLAR__procdff__DOLLAR__734__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[2] = __DOLLAR__procdff__DOLLAR__734__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[3] = __DOLLAR__procdff__DOLLAR__734__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[4] = __DOLLAR__procdff__DOLLAR__734__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[5] = __DOLLAR__procdff__DOLLAR__734__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[6] = __DOLLAR__procdff__DOLLAR__734__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[7] = __DOLLAR__procdff__DOLLAR__734__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[8] = __DOLLAR__procdff__DOLLAR__734__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__B[9] = __DOLLAR__procdff__DOLLAR__734__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[0] = __DOLLAR__procdff__DOLLAR__735__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[1] = __DOLLAR__procdff__DOLLAR__735__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[10] = __DOLLAR__procdff__DOLLAR__735__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[11] = __DOLLAR__procdff__DOLLAR__735__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[12] = __DOLLAR__procdff__DOLLAR__735__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[13] = __DOLLAR__procdff__DOLLAR__735__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[14] = __DOLLAR__procdff__DOLLAR__735__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[15] = __DOLLAR__procdff__DOLLAR__735__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[2] = __DOLLAR__procdff__DOLLAR__735__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[3] = __DOLLAR__procdff__DOLLAR__735__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[4] = __DOLLAR__procdff__DOLLAR__735__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[5] = __DOLLAR__procdff__DOLLAR__735__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[6] = __DOLLAR__procdff__DOLLAR__735__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[7] = __DOLLAR__procdff__DOLLAR__735__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[8] = __DOLLAR__procdff__DOLLAR__735__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__B[9] = __DOLLAR__procdff__DOLLAR__735__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[0] = __DOLLAR__procdff__DOLLAR__736__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[1] = __DOLLAR__procdff__DOLLAR__736__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[10] = __DOLLAR__procdff__DOLLAR__736__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[11] = __DOLLAR__procdff__DOLLAR__736__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[12] = __DOLLAR__procdff__DOLLAR__736__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[13] = __DOLLAR__procdff__DOLLAR__736__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[14] = __DOLLAR__procdff__DOLLAR__736__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[15] = __DOLLAR__procdff__DOLLAR__736__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[2] = __DOLLAR__procdff__DOLLAR__736__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[3] = __DOLLAR__procdff__DOLLAR__736__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[4] = __DOLLAR__procdff__DOLLAR__736__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[5] = __DOLLAR__procdff__DOLLAR__736__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[6] = __DOLLAR__procdff__DOLLAR__736__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[7] = __DOLLAR__procdff__DOLLAR__736__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[8] = __DOLLAR__procdff__DOLLAR__736__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__B[9] = __DOLLAR__procdff__DOLLAR__736__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[0] = __DOLLAR__procdff__DOLLAR__737__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[1] = __DOLLAR__procdff__DOLLAR__737__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[10] = __DOLLAR__procdff__DOLLAR__737__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[11] = __DOLLAR__procdff__DOLLAR__737__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[12] = __DOLLAR__procdff__DOLLAR__737__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[13] = __DOLLAR__procdff__DOLLAR__737__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[14] = __DOLLAR__procdff__DOLLAR__737__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[15] = __DOLLAR__procdff__DOLLAR__737__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[2] = __DOLLAR__procdff__DOLLAR__737__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[3] = __DOLLAR__procdff__DOLLAR__737__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[4] = __DOLLAR__procdff__DOLLAR__737__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[5] = __DOLLAR__procdff__DOLLAR__737__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[6] = __DOLLAR__procdff__DOLLAR__737__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[7] = __DOLLAR__procdff__DOLLAR__737__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[8] = __DOLLAR__procdff__DOLLAR__737__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__B[9] = __DOLLAR__procdff__DOLLAR__737__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[0] = __DOLLAR__procdff__DOLLAR__738__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[1] = __DOLLAR__procdff__DOLLAR__738__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[10] = __DOLLAR__procdff__DOLLAR__738__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[11] = __DOLLAR__procdff__DOLLAR__738__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[12] = __DOLLAR__procdff__DOLLAR__738__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[13] = __DOLLAR__procdff__DOLLAR__738__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[14] = __DOLLAR__procdff__DOLLAR__738__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[15] = __DOLLAR__procdff__DOLLAR__738__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[2] = __DOLLAR__procdff__DOLLAR__738__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[3] = __DOLLAR__procdff__DOLLAR__738__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[4] = __DOLLAR__procdff__DOLLAR__738__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[5] = __DOLLAR__procdff__DOLLAR__738__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[6] = __DOLLAR__procdff__DOLLAR__738__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[7] = __DOLLAR__procdff__DOLLAR__738__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[8] = __DOLLAR__procdff__DOLLAR__738__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__B[9] = __DOLLAR__procdff__DOLLAR__738__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[0] = __DOLLAR__procdff__DOLLAR__739__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[1] = __DOLLAR__procdff__DOLLAR__739__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[10] = __DOLLAR__procdff__DOLLAR__739__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[11] = __DOLLAR__procdff__DOLLAR__739__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[12] = __DOLLAR__procdff__DOLLAR__739__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[13] = __DOLLAR__procdff__DOLLAR__739__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[14] = __DOLLAR__procdff__DOLLAR__739__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[15] = __DOLLAR__procdff__DOLLAR__739__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[2] = __DOLLAR__procdff__DOLLAR__739__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[3] = __DOLLAR__procdff__DOLLAR__739__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[4] = __DOLLAR__procdff__DOLLAR__739__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[5] = __DOLLAR__procdff__DOLLAR__739__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[6] = __DOLLAR__procdff__DOLLAR__739__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[7] = __DOLLAR__procdff__DOLLAR__739__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[8] = __DOLLAR__procdff__DOLLAR__739__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__B[9] = __DOLLAR__procdff__DOLLAR__739__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[0] = __DOLLAR__procdff__DOLLAR__740__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[1] = __DOLLAR__procdff__DOLLAR__740__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[10] = __DOLLAR__procdff__DOLLAR__740__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[11] = __DOLLAR__procdff__DOLLAR__740__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[12] = __DOLLAR__procdff__DOLLAR__740__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[13] = __DOLLAR__procdff__DOLLAR__740__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[14] = __DOLLAR__procdff__DOLLAR__740__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[15] = __DOLLAR__procdff__DOLLAR__740__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[2] = __DOLLAR__procdff__DOLLAR__740__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[3] = __DOLLAR__procdff__DOLLAR__740__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[4] = __DOLLAR__procdff__DOLLAR__740__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[5] = __DOLLAR__procdff__DOLLAR__740__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[6] = __DOLLAR__procdff__DOLLAR__740__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[7] = __DOLLAR__procdff__DOLLAR__740__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[8] = __DOLLAR__procdff__DOLLAR__740__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__B[9] = __DOLLAR__procdff__DOLLAR__740__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[0] = __DOLLAR__procdff__DOLLAR__741__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[1] = __DOLLAR__procdff__DOLLAR__741__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[10] = __DOLLAR__procdff__DOLLAR__741__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[11] = __DOLLAR__procdff__DOLLAR__741__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[12] = __DOLLAR__procdff__DOLLAR__741__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[13] = __DOLLAR__procdff__DOLLAR__741__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[14] = __DOLLAR__procdff__DOLLAR__741__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[15] = __DOLLAR__procdff__DOLLAR__741__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[2] = __DOLLAR__procdff__DOLLAR__741__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[3] = __DOLLAR__procdff__DOLLAR__741__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[4] = __DOLLAR__procdff__DOLLAR__741__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[5] = __DOLLAR__procdff__DOLLAR__741__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[6] = __DOLLAR__procdff__DOLLAR__741__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[7] = __DOLLAR__procdff__DOLLAR__741__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[8] = __DOLLAR__procdff__DOLLAR__741__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__B[9] = __DOLLAR__procdff__DOLLAR__741__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[0] = __DOLLAR__procdff__DOLLAR__742__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[1] = __DOLLAR__procdff__DOLLAR__742__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[10] = __DOLLAR__procdff__DOLLAR__742__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[11] = __DOLLAR__procdff__DOLLAR__742__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[12] = __DOLLAR__procdff__DOLLAR__742__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[13] = __DOLLAR__procdff__DOLLAR__742__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[14] = __DOLLAR__procdff__DOLLAR__742__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[15] = __DOLLAR__procdff__DOLLAR__742__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[2] = __DOLLAR__procdff__DOLLAR__742__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[3] = __DOLLAR__procdff__DOLLAR__742__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[4] = __DOLLAR__procdff__DOLLAR__742__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[5] = __DOLLAR__procdff__DOLLAR__742__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[6] = __DOLLAR__procdff__DOLLAR__742__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[7] = __DOLLAR__procdff__DOLLAR__742__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[8] = __DOLLAR__procdff__DOLLAR__742__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__B[9] = __DOLLAR__procdff__DOLLAR__742__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[0] = __DOLLAR__procdff__DOLLAR__743__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[1] = __DOLLAR__procdff__DOLLAR__743__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[10] = __DOLLAR__procdff__DOLLAR__743__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[11] = __DOLLAR__procdff__DOLLAR__743__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[12] = __DOLLAR__procdff__DOLLAR__743__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[13] = __DOLLAR__procdff__DOLLAR__743__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[14] = __DOLLAR__procdff__DOLLAR__743__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[15] = __DOLLAR__procdff__DOLLAR__743__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[2] = __DOLLAR__procdff__DOLLAR__743__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[3] = __DOLLAR__procdff__DOLLAR__743__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[4] = __DOLLAR__procdff__DOLLAR__743__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[5] = __DOLLAR__procdff__DOLLAR__743__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[6] = __DOLLAR__procdff__DOLLAR__743__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[7] = __DOLLAR__procdff__DOLLAR__743__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[8] = __DOLLAR__procdff__DOLLAR__743__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__B[9] = __DOLLAR__procdff__DOLLAR__743__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[0] = __DOLLAR__procdff__DOLLAR__744__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[1] = __DOLLAR__procdff__DOLLAR__744__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[10] = __DOLLAR__procdff__DOLLAR__744__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[11] = __DOLLAR__procdff__DOLLAR__744__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[12] = __DOLLAR__procdff__DOLLAR__744__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[13] = __DOLLAR__procdff__DOLLAR__744__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[14] = __DOLLAR__procdff__DOLLAR__744__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[15] = __DOLLAR__procdff__DOLLAR__744__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[2] = __DOLLAR__procdff__DOLLAR__744__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[3] = __DOLLAR__procdff__DOLLAR__744__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[4] = __DOLLAR__procdff__DOLLAR__744__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[5] = __DOLLAR__procdff__DOLLAR__744__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[6] = __DOLLAR__procdff__DOLLAR__744__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[7] = __DOLLAR__procdff__DOLLAR__744__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[8] = __DOLLAR__procdff__DOLLAR__744__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__B[9] = __DOLLAR__procdff__DOLLAR__744__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[0] = __DOLLAR__procdff__DOLLAR__745__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[1] = __DOLLAR__procdff__DOLLAR__745__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[10] = __DOLLAR__procdff__DOLLAR__745__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[11] = __DOLLAR__procdff__DOLLAR__745__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[12] = __DOLLAR__procdff__DOLLAR__745__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[13] = __DOLLAR__procdff__DOLLAR__745__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[14] = __DOLLAR__procdff__DOLLAR__745__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[15] = __DOLLAR__procdff__DOLLAR__745__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[2] = __DOLLAR__procdff__DOLLAR__745__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[3] = __DOLLAR__procdff__DOLLAR__745__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[4] = __DOLLAR__procdff__DOLLAR__745__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[5] = __DOLLAR__procdff__DOLLAR__745__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[6] = __DOLLAR__procdff__DOLLAR__745__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[7] = __DOLLAR__procdff__DOLLAR__745__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[8] = __DOLLAR__procdff__DOLLAR__745__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__B[9] = __DOLLAR__procdff__DOLLAR__745__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[0] = __DOLLAR__procdff__DOLLAR__746__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[1] = __DOLLAR__procdff__DOLLAR__746__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[10] = __DOLLAR__procdff__DOLLAR__746__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[11] = __DOLLAR__procdff__DOLLAR__746__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[12] = __DOLLAR__procdff__DOLLAR__746__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[13] = __DOLLAR__procdff__DOLLAR__746__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[14] = __DOLLAR__procdff__DOLLAR__746__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[15] = __DOLLAR__procdff__DOLLAR__746__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[2] = __DOLLAR__procdff__DOLLAR__746__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[3] = __DOLLAR__procdff__DOLLAR__746__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[4] = __DOLLAR__procdff__DOLLAR__746__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[5] = __DOLLAR__procdff__DOLLAR__746__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[6] = __DOLLAR__procdff__DOLLAR__746__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[7] = __DOLLAR__procdff__DOLLAR__746__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[8] = __DOLLAR__procdff__DOLLAR__746__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__B[9] = __DOLLAR__procdff__DOLLAR__746__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[0] = __DOLLAR__procdff__DOLLAR__747__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[1] = __DOLLAR__procdff__DOLLAR__747__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[10] = __DOLLAR__procdff__DOLLAR__747__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[11] = __DOLLAR__procdff__DOLLAR__747__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[12] = __DOLLAR__procdff__DOLLAR__747__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[13] = __DOLLAR__procdff__DOLLAR__747__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[14] = __DOLLAR__procdff__DOLLAR__747__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[15] = __DOLLAR__procdff__DOLLAR__747__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[2] = __DOLLAR__procdff__DOLLAR__747__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[3] = __DOLLAR__procdff__DOLLAR__747__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[4] = __DOLLAR__procdff__DOLLAR__747__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[5] = __DOLLAR__procdff__DOLLAR__747__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[6] = __DOLLAR__procdff__DOLLAR__747__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[7] = __DOLLAR__procdff__DOLLAR__747__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[8] = __DOLLAR__procdff__DOLLAR__747__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__B[9] = __DOLLAR__procdff__DOLLAR__747__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[0] = __DOLLAR__procdff__DOLLAR__748__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[1] = __DOLLAR__procdff__DOLLAR__748__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[10] = __DOLLAR__procdff__DOLLAR__748__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[11] = __DOLLAR__procdff__DOLLAR__748__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[12] = __DOLLAR__procdff__DOLLAR__748__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[13] = __DOLLAR__procdff__DOLLAR__748__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[14] = __DOLLAR__procdff__DOLLAR__748__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[15] = __DOLLAR__procdff__DOLLAR__748__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[2] = __DOLLAR__procdff__DOLLAR__748__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[3] = __DOLLAR__procdff__DOLLAR__748__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[4] = __DOLLAR__procdff__DOLLAR__748__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[5] = __DOLLAR__procdff__DOLLAR__748__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[6] = __DOLLAR__procdff__DOLLAR__748__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[7] = __DOLLAR__procdff__DOLLAR__748__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[8] = __DOLLAR__procdff__DOLLAR__748__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__B[9] = __DOLLAR__procdff__DOLLAR__748__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[0] = __DOLLAR__procdff__DOLLAR__749__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[1] = __DOLLAR__procdff__DOLLAR__749__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[10] = __DOLLAR__procdff__DOLLAR__749__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[11] = __DOLLAR__procdff__DOLLAR__749__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[12] = __DOLLAR__procdff__DOLLAR__749__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[13] = __DOLLAR__procdff__DOLLAR__749__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[14] = __DOLLAR__procdff__DOLLAR__749__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[15] = __DOLLAR__procdff__DOLLAR__749__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[2] = __DOLLAR__procdff__DOLLAR__749__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[3] = __DOLLAR__procdff__DOLLAR__749__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[4] = __DOLLAR__procdff__DOLLAR__749__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[5] = __DOLLAR__procdff__DOLLAR__749__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[6] = __DOLLAR__procdff__DOLLAR__749__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[7] = __DOLLAR__procdff__DOLLAR__749__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[8] = __DOLLAR__procdff__DOLLAR__749__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__B[9] = __DOLLAR__procdff__DOLLAR__749__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[0] = __DOLLAR__procdff__DOLLAR__750__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[1] = __DOLLAR__procdff__DOLLAR__750__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[10] = __DOLLAR__procdff__DOLLAR__750__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[11] = __DOLLAR__procdff__DOLLAR__750__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[12] = __DOLLAR__procdff__DOLLAR__750__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[13] = __DOLLAR__procdff__DOLLAR__750__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[14] = __DOLLAR__procdff__DOLLAR__750__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[15] = __DOLLAR__procdff__DOLLAR__750__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[2] = __DOLLAR__procdff__DOLLAR__750__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[3] = __DOLLAR__procdff__DOLLAR__750__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[4] = __DOLLAR__procdff__DOLLAR__750__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[5] = __DOLLAR__procdff__DOLLAR__750__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[6] = __DOLLAR__procdff__DOLLAR__750__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[7] = __DOLLAR__procdff__DOLLAR__750__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[8] = __DOLLAR__procdff__DOLLAR__750__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__B[9] = __DOLLAR__procdff__DOLLAR__750__Q[9];
  assign __DOLLAR__procdff__DOLLAR__751__D[0] = __DOLLAR__procmux__DOLLAR__522__Y[0];
  assign __DOLLAR__procdff__DOLLAR__751__D[1] = __DOLLAR__procmux__DOLLAR__522__Y[1];
  assign __DOLLAR__procdff__DOLLAR__751__D[10] = __DOLLAR__procmux__DOLLAR__522__Y[10];
  assign __DOLLAR__procdff__DOLLAR__751__D[11] = __DOLLAR__procmux__DOLLAR__522__Y[11];
  assign __DOLLAR__procdff__DOLLAR__751__D[12] = __DOLLAR__procmux__DOLLAR__522__Y[12];
  assign __DOLLAR__procdff__DOLLAR__751__D[13] = __DOLLAR__procmux__DOLLAR__522__Y[13];
  assign __DOLLAR__procdff__DOLLAR__751__D[14] = __DOLLAR__procmux__DOLLAR__522__Y[14];
  assign __DOLLAR__procdff__DOLLAR__751__D[15] = __DOLLAR__procmux__DOLLAR__522__Y[15];
  assign __DOLLAR__procdff__DOLLAR__751__D[16] = __DOLLAR__procmux__DOLLAR__522__Y[16];
  assign __DOLLAR__procdff__DOLLAR__751__D[17] = __DOLLAR__procmux__DOLLAR__522__Y[17];
  assign __DOLLAR__procdff__DOLLAR__751__D[18] = __DOLLAR__procmux__DOLLAR__522__Y[18];
  assign __DOLLAR__procdff__DOLLAR__751__D[19] = __DOLLAR__procmux__DOLLAR__522__Y[19];
  assign __DOLLAR__procdff__DOLLAR__751__D[2] = __DOLLAR__procmux__DOLLAR__522__Y[2];
  assign __DOLLAR__procdff__DOLLAR__751__D[20] = __DOLLAR__procmux__DOLLAR__522__Y[20];
  assign __DOLLAR__procdff__DOLLAR__751__D[21] = __DOLLAR__procmux__DOLLAR__522__Y[21];
  assign __DOLLAR__procdff__DOLLAR__751__D[22] = __DOLLAR__procmux__DOLLAR__522__Y[22];
  assign __DOLLAR__procdff__DOLLAR__751__D[23] = __DOLLAR__procmux__DOLLAR__522__Y[23];
  assign __DOLLAR__procdff__DOLLAR__751__D[24] = __DOLLAR__procmux__DOLLAR__522__Y[24];
  assign __DOLLAR__procdff__DOLLAR__751__D[25] = __DOLLAR__procmux__DOLLAR__522__Y[25];
  assign __DOLLAR__procdff__DOLLAR__751__D[26] = __DOLLAR__procmux__DOLLAR__522__Y[26];
  assign __DOLLAR__procdff__DOLLAR__751__D[27] = __DOLLAR__procmux__DOLLAR__522__Y[27];
  assign __DOLLAR__procdff__DOLLAR__751__D[28] = __DOLLAR__procmux__DOLLAR__522__Y[28];
  assign __DOLLAR__procdff__DOLLAR__751__D[29] = __DOLLAR__procmux__DOLLAR__522__Y[29];
  assign __DOLLAR__procdff__DOLLAR__751__D[3] = __DOLLAR__procmux__DOLLAR__522__Y[3];
  assign __DOLLAR__procdff__DOLLAR__751__D[30] = __DOLLAR__procmux__DOLLAR__522__Y[30];
  assign __DOLLAR__procdff__DOLLAR__751__D[31] = __DOLLAR__procmux__DOLLAR__522__Y[31];
  assign __DOLLAR__procdff__DOLLAR__751__D[32] = __DOLLAR__procmux__DOLLAR__515__Y[0];
  assign __DOLLAR__procdff__DOLLAR__751__D[33] = __DOLLAR__procmux__DOLLAR__515__Y[1];
  assign __DOLLAR__procdff__DOLLAR__751__D[34] = __DOLLAR__procmux__DOLLAR__515__Y[2];
  assign __DOLLAR__procdff__DOLLAR__751__D[35] = __DOLLAR__procmux__DOLLAR__515__Y[3];
  assign __DOLLAR__procdff__DOLLAR__751__D[36] = __DOLLAR__procmux__DOLLAR__515__Y[4];
  assign __DOLLAR__procdff__DOLLAR__751__D[37] = __DOLLAR__procmux__DOLLAR__515__Y[5];
  assign __DOLLAR__procdff__DOLLAR__751__D[38] = __DOLLAR__procmux__DOLLAR__515__Y[6];
  assign __DOLLAR__procdff__DOLLAR__751__D[39] = __DOLLAR__procmux__DOLLAR__515__Y[7];
  assign __DOLLAR__procdff__DOLLAR__751__D[4] = __DOLLAR__procmux__DOLLAR__522__Y[4];
  assign __DOLLAR__procdff__DOLLAR__751__D[40] = __DOLLAR__procmux__DOLLAR__515__Y[8];
  assign __DOLLAR__procdff__DOLLAR__751__D[41] = __DOLLAR__procmux__DOLLAR__515__Y[9];
  assign __DOLLAR__procdff__DOLLAR__751__D[42] = __DOLLAR__procmux__DOLLAR__515__Y[10];
  assign __DOLLAR__procdff__DOLLAR__751__D[43] = __DOLLAR__procmux__DOLLAR__515__Y[11];
  assign __DOLLAR__procdff__DOLLAR__751__D[44] = __DOLLAR__procmux__DOLLAR__515__Y[12];
  assign __DOLLAR__procdff__DOLLAR__751__D[45] = __DOLLAR__procmux__DOLLAR__515__Y[13];
  assign __DOLLAR__procdff__DOLLAR__751__D[46] = __DOLLAR__procmux__DOLLAR__515__Y[14];
  assign __DOLLAR__procdff__DOLLAR__751__D[47] = __DOLLAR__procmux__DOLLAR__515__Y[15];
  assign __DOLLAR__procdff__DOLLAR__751__D[48] = __DOLLAR__procmux__DOLLAR__515__Y[16];
  assign __DOLLAR__procdff__DOLLAR__751__D[49] = __DOLLAR__procmux__DOLLAR__515__Y[17];
  assign __DOLLAR__procdff__DOLLAR__751__D[5] = __DOLLAR__procmux__DOLLAR__522__Y[5];
  assign __DOLLAR__procdff__DOLLAR__751__D[50] = __DOLLAR__procmux__DOLLAR__515__Y[18];
  assign __DOLLAR__procdff__DOLLAR__751__D[51] = __DOLLAR__procmux__DOLLAR__515__Y[19];
  assign __DOLLAR__procdff__DOLLAR__751__D[52] = __DOLLAR__procmux__DOLLAR__515__Y[20];
  assign __DOLLAR__procdff__DOLLAR__751__D[53] = __DOLLAR__procmux__DOLLAR__515__Y[21];
  assign __DOLLAR__procdff__DOLLAR__751__D[54] = __DOLLAR__procmux__DOLLAR__515__Y[22];
  assign __DOLLAR__procdff__DOLLAR__751__D[55] = __DOLLAR__procmux__DOLLAR__515__Y[23];
  assign __DOLLAR__procdff__DOLLAR__751__D[56] = __DOLLAR__procmux__DOLLAR__515__Y[24];
  assign __DOLLAR__procdff__DOLLAR__751__D[57] = __DOLLAR__procmux__DOLLAR__515__Y[25];
  assign __DOLLAR__procdff__DOLLAR__751__D[58] = __DOLLAR__procmux__DOLLAR__515__Y[26];
  assign __DOLLAR__procdff__DOLLAR__751__D[59] = __DOLLAR__procmux__DOLLAR__515__Y[27];
  assign __DOLLAR__procdff__DOLLAR__751__D[6] = __DOLLAR__procmux__DOLLAR__522__Y[6];
  assign __DOLLAR__procdff__DOLLAR__751__D[60] = __DOLLAR__procmux__DOLLAR__515__Y[28];
  assign __DOLLAR__procdff__DOLLAR__751__D[61] = __DOLLAR__procmux__DOLLAR__515__Y[29];
  assign __DOLLAR__procdff__DOLLAR__751__D[62] = __DOLLAR__procmux__DOLLAR__515__Y[30];
  assign __DOLLAR__procdff__DOLLAR__751__D[63] = __DOLLAR__procmux__DOLLAR__515__Y[31];
  assign __DOLLAR__procdff__DOLLAR__751__D[7] = __DOLLAR__procmux__DOLLAR__522__Y[7];
  assign __DOLLAR__procdff__DOLLAR__751__D[8] = __DOLLAR__procmux__DOLLAR__522__Y[8];
  assign __DOLLAR__procdff__DOLLAR__751__D[9] = __DOLLAR__procmux__DOLLAR__522__Y[9];
  assign __DOLLAR__procmux__DOLLAR__507_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__508_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__509_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__510_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__520__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__522__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign config_sb_res[0] = __DOLLAR__procdff__DOLLAR__751__Q[0];
  assign __DOLLAR__procmux__DOLLAR__507_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__508_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__509_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__510_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__520__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__522__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign config_sb_res[1] = __DOLLAR__procdff__DOLLAR__751__Q[1];
  assign __DOLLAR__procmux__DOLLAR__482_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__483_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__484_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__485_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__520__A[10] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__522__A[10] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign config_sb_res[10] = __DOLLAR__procdff__DOLLAR__751__Q[10];
  assign __DOLLAR__procmux__DOLLAR__482_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__483_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__484_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__485_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__520__A[11] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__522__A[11] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign config_sb_res[11] = __DOLLAR__procdff__DOLLAR__751__Q[11];
  assign __DOLLAR__procmux__DOLLAR__477_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__478_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__479_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__480_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__520__A[12] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__522__A[12] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign config_sb_res[12] = __DOLLAR__procdff__DOLLAR__751__Q[12];
  assign __DOLLAR__procmux__DOLLAR__477_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__478_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__479_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__480_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__520__A[13] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__522__A[13] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign config_sb_res[13] = __DOLLAR__procdff__DOLLAR__751__Q[13];
  assign __DOLLAR__procmux__DOLLAR__472_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__473_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__474_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__475_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__520__A[14] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__522__A[14] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign config_sb_res[14] = __DOLLAR__procdff__DOLLAR__751__Q[14];
  assign __DOLLAR__procmux__DOLLAR__472_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__473_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__474_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__475_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__520__A[15] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__522__A[15] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign config_sb_res[15] = __DOLLAR__procdff__DOLLAR__751__Q[15];
  assign __DOLLAR__procmux__DOLLAR__467_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__468_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__469_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__470_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__520__A[16] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__522__A[16] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign config_sb_res[16] = __DOLLAR__procdff__DOLLAR__751__Q[16];
  assign __DOLLAR__procmux__DOLLAR__467_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__468_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__469_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__470_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__520__A[17] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__522__A[17] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign config_sb_res[17] = __DOLLAR__procdff__DOLLAR__751__Q[17];
  assign __DOLLAR__procmux__DOLLAR__462_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__463_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__464_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__465_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__520__A[18] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__522__A[18] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign config_sb_res[18] = __DOLLAR__procdff__DOLLAR__751__Q[18];
  assign __DOLLAR__procmux__DOLLAR__462_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__463_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__464_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__465_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__520__A[19] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__522__A[19] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign config_sb_res[19] = __DOLLAR__procdff__DOLLAR__751__Q[19];
  assign __DOLLAR__procmux__DOLLAR__502_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__503_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__504_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__505_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__520__A[2] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__522__A[2] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign config_sb_res[2] = __DOLLAR__procdff__DOLLAR__751__Q[2];
  assign __DOLLAR__procmux__DOLLAR__457_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__458_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__459_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__460_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__520__A[20] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__522__A[20] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign config_sb_res[20] = __DOLLAR__procdff__DOLLAR__751__Q[20];
  assign __DOLLAR__procmux__DOLLAR__457_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__458_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__459_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__460_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__520__A[21] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__522__A[21] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign config_sb_res[21] = __DOLLAR__procdff__DOLLAR__751__Q[21];
  assign __DOLLAR__procmux__DOLLAR__452_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__453_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__454_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__455_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__520__A[22] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__522__A[22] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign config_sb_res[22] = __DOLLAR__procdff__DOLLAR__751__Q[22];
  assign __DOLLAR__procmux__DOLLAR__452_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__453_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__454_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__455_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__520__A[23] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__522__A[23] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign config_sb_res[23] = __DOLLAR__procdff__DOLLAR__751__Q[23];
  assign __DOLLAR__procmux__DOLLAR__447_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__448_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__449_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__450_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__520__A[24] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__522__A[24] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign config_sb_res[24] = __DOLLAR__procdff__DOLLAR__751__Q[24];
  assign __DOLLAR__procmux__DOLLAR__447_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__448_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__449_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__450_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__520__A[25] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__522__A[25] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign config_sb_res[25] = __DOLLAR__procdff__DOLLAR__751__Q[25];
  assign __DOLLAR__procmux__DOLLAR__442_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__443_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__444_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__445_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__520__A[26] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__522__A[26] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign config_sb_res[26] = __DOLLAR__procdff__DOLLAR__751__Q[26];
  assign __DOLLAR__procmux__DOLLAR__442_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__443_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__444_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__445_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__520__A[27] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__522__A[27] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign config_sb_res[27] = __DOLLAR__procdff__DOLLAR__751__Q[27];
  assign __DOLLAR__procmux__DOLLAR__437_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__438_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__439_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__440_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__520__A[28] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__522__A[28] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign config_sb_res[28] = __DOLLAR__procdff__DOLLAR__751__Q[28];
  assign __DOLLAR__procmux__DOLLAR__437_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__438_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__439_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__440_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__520__A[29] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__522__A[29] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign config_sb_res[29] = __DOLLAR__procdff__DOLLAR__751__Q[29];
  assign __DOLLAR__procmux__DOLLAR__502_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__503_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__504_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__505_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__520__A[3] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__522__A[3] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign config_sb_res[3] = __DOLLAR__procdff__DOLLAR__751__Q[3];
  assign __DOLLAR__procmux__DOLLAR__432_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__433_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__434_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__435_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__520__A[30] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__522__A[30] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign config_sb_res[30] = __DOLLAR__procdff__DOLLAR__751__Q[30];
  assign __DOLLAR__procmux__DOLLAR__432_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__433_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__434_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__435_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__520__A[31] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__522__A[31] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign config_sb_res[31] = __DOLLAR__procdff__DOLLAR__751__Q[31];
  assign __DOLLAR__procmux__DOLLAR__427_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__428_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__429_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__430_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__513__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__515__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign config_sb_res[32] = __DOLLAR__procdff__DOLLAR__751__Q[32];
  assign __DOLLAR__procmux__DOLLAR__427_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__428_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__429_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__430_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__513__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__515__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign config_sb_res[33] = __DOLLAR__procdff__DOLLAR__751__Q[33];
  assign __DOLLAR__procmux__DOLLAR__422_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__423_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__424_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__425_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__513__A[2] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__515__A[2] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign config_sb_res[34] = __DOLLAR__procdff__DOLLAR__751__Q[34];
  assign __DOLLAR__procmux__DOLLAR__422_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__423_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__424_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__425_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__513__A[3] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__515__A[3] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign config_sb_res[35] = __DOLLAR__procdff__DOLLAR__751__Q[35];
  assign __DOLLAR__procmux__DOLLAR__417_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__418_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__419_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__420_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__513__A[4] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__515__A[4] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign config_sb_res[36] = __DOLLAR__procdff__DOLLAR__751__Q[36];
  assign __DOLLAR__procmux__DOLLAR__417_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__418_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__419_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__420_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__513__A[5] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__515__A[5] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign config_sb_res[37] = __DOLLAR__procdff__DOLLAR__751__Q[37];
  assign __DOLLAR__procmux__DOLLAR__412_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__413_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__414_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__415_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__513__A[6] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__515__A[6] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign config_sb_res[38] = __DOLLAR__procdff__DOLLAR__751__Q[38];
  assign __DOLLAR__procmux__DOLLAR__412_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__413_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__414_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__415_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__513__A[7] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__515__A[7] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign config_sb_res[39] = __DOLLAR__procdff__DOLLAR__751__Q[39];
  assign __DOLLAR__procmux__DOLLAR__497_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__498_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__499_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__500_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__520__A[4] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__522__A[4] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign config_sb_res[4] = __DOLLAR__procdff__DOLLAR__751__Q[4];
  assign __DOLLAR__procmux__DOLLAR__513__A[8] = __DOLLAR__procdff__DOLLAR__751__Q[40];
  assign __DOLLAR__procmux__DOLLAR__515__A[8] = __DOLLAR__procdff__DOLLAR__751__Q[40];
  assign config_sb_res[40] = __DOLLAR__procdff__DOLLAR__751__Q[40];
  assign __DOLLAR__procmux__DOLLAR__513__A[9] = __DOLLAR__procdff__DOLLAR__751__Q[41];
  assign __DOLLAR__procmux__DOLLAR__515__A[9] = __DOLLAR__procdff__DOLLAR__751__Q[41];
  assign config_sb_res[41] = __DOLLAR__procdff__DOLLAR__751__Q[41];
  assign __DOLLAR__procmux__DOLLAR__513__A[10] = __DOLLAR__procdff__DOLLAR__751__Q[42];
  assign __DOLLAR__procmux__DOLLAR__515__A[10] = __DOLLAR__procdff__DOLLAR__751__Q[42];
  assign config_sb_res[42] = __DOLLAR__procdff__DOLLAR__751__Q[42];
  assign __DOLLAR__procmux__DOLLAR__513__A[11] = __DOLLAR__procdff__DOLLAR__751__Q[43];
  assign __DOLLAR__procmux__DOLLAR__515__A[11] = __DOLLAR__procdff__DOLLAR__751__Q[43];
  assign config_sb_res[43] = __DOLLAR__procdff__DOLLAR__751__Q[43];
  assign __DOLLAR__procmux__DOLLAR__513__A[12] = __DOLLAR__procdff__DOLLAR__751__Q[44];
  assign __DOLLAR__procmux__DOLLAR__515__A[12] = __DOLLAR__procdff__DOLLAR__751__Q[44];
  assign config_sb_res[44] = __DOLLAR__procdff__DOLLAR__751__Q[44];
  assign __DOLLAR__procmux__DOLLAR__513__A[13] = __DOLLAR__procdff__DOLLAR__751__Q[45];
  assign __DOLLAR__procmux__DOLLAR__515__A[13] = __DOLLAR__procdff__DOLLAR__751__Q[45];
  assign config_sb_res[45] = __DOLLAR__procdff__DOLLAR__751__Q[45];
  assign __DOLLAR__procmux__DOLLAR__513__A[14] = __DOLLAR__procdff__DOLLAR__751__Q[46];
  assign __DOLLAR__procmux__DOLLAR__515__A[14] = __DOLLAR__procdff__DOLLAR__751__Q[46];
  assign config_sb_res[46] = __DOLLAR__procdff__DOLLAR__751__Q[46];
  assign __DOLLAR__procmux__DOLLAR__513__A[15] = __DOLLAR__procdff__DOLLAR__751__Q[47];
  assign __DOLLAR__procmux__DOLLAR__515__A[15] = __DOLLAR__procdff__DOLLAR__751__Q[47];
  assign config_sb_res[47] = __DOLLAR__procdff__DOLLAR__751__Q[47];
  assign __DOLLAR__procmux__DOLLAR__513__A[16] = __DOLLAR__procdff__DOLLAR__751__Q[48];
  assign __DOLLAR__procmux__DOLLAR__515__A[16] = __DOLLAR__procdff__DOLLAR__751__Q[48];
  assign config_sb_res[48] = __DOLLAR__procdff__DOLLAR__751__Q[48];
  assign __DOLLAR__procmux__DOLLAR__513__A[17] = __DOLLAR__procdff__DOLLAR__751__Q[49];
  assign __DOLLAR__procmux__DOLLAR__515__A[17] = __DOLLAR__procdff__DOLLAR__751__Q[49];
  assign config_sb_res[49] = __DOLLAR__procdff__DOLLAR__751__Q[49];
  assign __DOLLAR__procmux__DOLLAR__497_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__498_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__499_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__500_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__520__A[5] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__522__A[5] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign config_sb_res[5] = __DOLLAR__procdff__DOLLAR__751__Q[5];
  assign __DOLLAR__procmux__DOLLAR__513__A[18] = __DOLLAR__procdff__DOLLAR__751__Q[50];
  assign __DOLLAR__procmux__DOLLAR__515__A[18] = __DOLLAR__procdff__DOLLAR__751__Q[50];
  assign config_sb_res[50] = __DOLLAR__procdff__DOLLAR__751__Q[50];
  assign __DOLLAR__procmux__DOLLAR__513__A[19] = __DOLLAR__procdff__DOLLAR__751__Q[51];
  assign __DOLLAR__procmux__DOLLAR__515__A[19] = __DOLLAR__procdff__DOLLAR__751__Q[51];
  assign config_sb_res[51] = __DOLLAR__procdff__DOLLAR__751__Q[51];
  assign __DOLLAR__procmux__DOLLAR__513__A[20] = __DOLLAR__procdff__DOLLAR__751__Q[52];
  assign __DOLLAR__procmux__DOLLAR__515__A[20] = __DOLLAR__procdff__DOLLAR__751__Q[52];
  assign config_sb_res[52] = __DOLLAR__procdff__DOLLAR__751__Q[52];
  assign __DOLLAR__procmux__DOLLAR__513__A[21] = __DOLLAR__procdff__DOLLAR__751__Q[53];
  assign __DOLLAR__procmux__DOLLAR__515__A[21] = __DOLLAR__procdff__DOLLAR__751__Q[53];
  assign config_sb_res[53] = __DOLLAR__procdff__DOLLAR__751__Q[53];
  assign __DOLLAR__procmux__DOLLAR__513__A[22] = __DOLLAR__procdff__DOLLAR__751__Q[54];
  assign __DOLLAR__procmux__DOLLAR__515__A[22] = __DOLLAR__procdff__DOLLAR__751__Q[54];
  assign config_sb_res[54] = __DOLLAR__procdff__DOLLAR__751__Q[54];
  assign __DOLLAR__procmux__DOLLAR__513__A[23] = __DOLLAR__procdff__DOLLAR__751__Q[55];
  assign __DOLLAR__procmux__DOLLAR__515__A[23] = __DOLLAR__procdff__DOLLAR__751__Q[55];
  assign config_sb_res[55] = __DOLLAR__procdff__DOLLAR__751__Q[55];
  assign __DOLLAR__procmux__DOLLAR__513__A[24] = __DOLLAR__procdff__DOLLAR__751__Q[56];
  assign __DOLLAR__procmux__DOLLAR__515__A[24] = __DOLLAR__procdff__DOLLAR__751__Q[56];
  assign config_sb_res[56] = __DOLLAR__procdff__DOLLAR__751__Q[56];
  assign __DOLLAR__procmux__DOLLAR__513__A[25] = __DOLLAR__procdff__DOLLAR__751__Q[57];
  assign __DOLLAR__procmux__DOLLAR__515__A[25] = __DOLLAR__procdff__DOLLAR__751__Q[57];
  assign config_sb_res[57] = __DOLLAR__procdff__DOLLAR__751__Q[57];
  assign __DOLLAR__procmux__DOLLAR__513__A[26] = __DOLLAR__procdff__DOLLAR__751__Q[58];
  assign __DOLLAR__procmux__DOLLAR__515__A[26] = __DOLLAR__procdff__DOLLAR__751__Q[58];
  assign config_sb_res[58] = __DOLLAR__procdff__DOLLAR__751__Q[58];
  assign __DOLLAR__procmux__DOLLAR__513__A[27] = __DOLLAR__procdff__DOLLAR__751__Q[59];
  assign __DOLLAR__procmux__DOLLAR__515__A[27] = __DOLLAR__procdff__DOLLAR__751__Q[59];
  assign config_sb_res[59] = __DOLLAR__procdff__DOLLAR__751__Q[59];
  assign __DOLLAR__procmux__DOLLAR__492_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__493_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__494_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__495_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__520__A[6] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__522__A[6] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign config_sb_res[6] = __DOLLAR__procdff__DOLLAR__751__Q[6];
  assign __DOLLAR__procmux__DOLLAR__513__A[28] = __DOLLAR__procdff__DOLLAR__751__Q[60];
  assign __DOLLAR__procmux__DOLLAR__515__A[28] = __DOLLAR__procdff__DOLLAR__751__Q[60];
  assign config_sb_res[60] = __DOLLAR__procdff__DOLLAR__751__Q[60];
  assign __DOLLAR__procmux__DOLLAR__513__A[29] = __DOLLAR__procdff__DOLLAR__751__Q[61];
  assign __DOLLAR__procmux__DOLLAR__515__A[29] = __DOLLAR__procdff__DOLLAR__751__Q[61];
  assign config_sb_res[61] = __DOLLAR__procdff__DOLLAR__751__Q[61];
  assign __DOLLAR__procmux__DOLLAR__513__A[30] = __DOLLAR__procdff__DOLLAR__751__Q[62];
  assign __DOLLAR__procmux__DOLLAR__515__A[30] = __DOLLAR__procdff__DOLLAR__751__Q[62];
  assign config_sb_res[62] = __DOLLAR__procdff__DOLLAR__751__Q[62];
  assign __DOLLAR__procmux__DOLLAR__513__A[31] = __DOLLAR__procdff__DOLLAR__751__Q[63];
  assign __DOLLAR__procmux__DOLLAR__515__A[31] = __DOLLAR__procdff__DOLLAR__751__Q[63];
  assign config_sb_res[63] = __DOLLAR__procdff__DOLLAR__751__Q[63];
  assign __DOLLAR__procmux__DOLLAR__492_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__493_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__494_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__495_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__520__A[7] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__522__A[7] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign config_sb_res[7] = __DOLLAR__procdff__DOLLAR__751__Q[7];
  assign __DOLLAR__procmux__DOLLAR__487_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__488_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__489_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__490_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__520__A[8] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__522__A[8] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign config_sb_res[8] = __DOLLAR__procdff__DOLLAR__751__Q[8];
  assign __DOLLAR__procmux__DOLLAR__487_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__488_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__489_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__490_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__520__A[9] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__522__A[9] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign config_sb_res[9] = __DOLLAR__procdff__DOLLAR__751__Q[9];
  assign __DOLLAR__procmux__DOLLAR__513__B[0] = config_data[0];
  assign __DOLLAR__procmux__DOLLAR__513__B[1] = config_data[1];
  assign __DOLLAR__procmux__DOLLAR__513__B[10] = config_data[10];
  assign __DOLLAR__procmux__DOLLAR__513__B[11] = config_data[11];
  assign __DOLLAR__procmux__DOLLAR__513__B[12] = config_data[12];
  assign __DOLLAR__procmux__DOLLAR__513__B[13] = config_data[13];
  assign __DOLLAR__procmux__DOLLAR__513__B[14] = config_data[14];
  assign __DOLLAR__procmux__DOLLAR__513__B[15] = config_data[15];
  assign __DOLLAR__procmux__DOLLAR__513__B[16] = config_data[16];
  assign __DOLLAR__procmux__DOLLAR__513__B[17] = config_data[17];
  assign __DOLLAR__procmux__DOLLAR__513__B[18] = config_data[18];
  assign __DOLLAR__procmux__DOLLAR__513__B[19] = config_data[19];
  assign __DOLLAR__procmux__DOLLAR__513__B[2] = config_data[2];
  assign __DOLLAR__procmux__DOLLAR__513__B[20] = config_data[20];
  assign __DOLLAR__procmux__DOLLAR__513__B[21] = config_data[21];
  assign __DOLLAR__procmux__DOLLAR__513__B[22] = config_data[22];
  assign __DOLLAR__procmux__DOLLAR__513__B[23] = config_data[23];
  assign __DOLLAR__procmux__DOLLAR__513__B[24] = config_data[24];
  assign __DOLLAR__procmux__DOLLAR__513__B[25] = config_data[25];
  assign __DOLLAR__procmux__DOLLAR__513__B[26] = config_data[26];
  assign __DOLLAR__procmux__DOLLAR__513__B[27] = config_data[27];
  assign __DOLLAR__procmux__DOLLAR__513__B[28] = config_data[28];
  assign __DOLLAR__procmux__DOLLAR__513__B[29] = config_data[29];
  assign __DOLLAR__procmux__DOLLAR__513__B[3] = config_data[3];
  assign __DOLLAR__procmux__DOLLAR__513__B[30] = config_data[30];
  assign __DOLLAR__procmux__DOLLAR__513__B[31] = config_data[31];
  assign __DOLLAR__procmux__DOLLAR__513__B[4] = config_data[4];
  assign __DOLLAR__procmux__DOLLAR__513__B[5] = config_data[5];
  assign __DOLLAR__procmux__DOLLAR__513__B[6] = config_data[6];
  assign __DOLLAR__procmux__DOLLAR__513__B[7] = config_data[7];
  assign __DOLLAR__procmux__DOLLAR__513__B[8] = config_data[8];
  assign __DOLLAR__procmux__DOLLAR__513__B[9] = config_data[9];
  assign __DOLLAR__procmux__DOLLAR__515__B[0] = __DOLLAR__procmux__DOLLAR__513__Y[0];
  assign __DOLLAR__procmux__DOLLAR__515__B[1] = __DOLLAR__procmux__DOLLAR__513__Y[1];
  assign __DOLLAR__procmux__DOLLAR__515__B[10] = __DOLLAR__procmux__DOLLAR__513__Y[10];
  assign __DOLLAR__procmux__DOLLAR__515__B[11] = __DOLLAR__procmux__DOLLAR__513__Y[11];
  assign __DOLLAR__procmux__DOLLAR__515__B[12] = __DOLLAR__procmux__DOLLAR__513__Y[12];
  assign __DOLLAR__procmux__DOLLAR__515__B[13] = __DOLLAR__procmux__DOLLAR__513__Y[13];
  assign __DOLLAR__procmux__DOLLAR__515__B[14] = __DOLLAR__procmux__DOLLAR__513__Y[14];
  assign __DOLLAR__procmux__DOLLAR__515__B[15] = __DOLLAR__procmux__DOLLAR__513__Y[15];
  assign __DOLLAR__procmux__DOLLAR__515__B[16] = __DOLLAR__procmux__DOLLAR__513__Y[16];
  assign __DOLLAR__procmux__DOLLAR__515__B[17] = __DOLLAR__procmux__DOLLAR__513__Y[17];
  assign __DOLLAR__procmux__DOLLAR__515__B[18] = __DOLLAR__procmux__DOLLAR__513__Y[18];
  assign __DOLLAR__procmux__DOLLAR__515__B[19] = __DOLLAR__procmux__DOLLAR__513__Y[19];
  assign __DOLLAR__procmux__DOLLAR__515__B[2] = __DOLLAR__procmux__DOLLAR__513__Y[2];
  assign __DOLLAR__procmux__DOLLAR__515__B[20] = __DOLLAR__procmux__DOLLAR__513__Y[20];
  assign __DOLLAR__procmux__DOLLAR__515__B[21] = __DOLLAR__procmux__DOLLAR__513__Y[21];
  assign __DOLLAR__procmux__DOLLAR__515__B[22] = __DOLLAR__procmux__DOLLAR__513__Y[22];
  assign __DOLLAR__procmux__DOLLAR__515__B[23] = __DOLLAR__procmux__DOLLAR__513__Y[23];
  assign __DOLLAR__procmux__DOLLAR__515__B[24] = __DOLLAR__procmux__DOLLAR__513__Y[24];
  assign __DOLLAR__procmux__DOLLAR__515__B[25] = __DOLLAR__procmux__DOLLAR__513__Y[25];
  assign __DOLLAR__procmux__DOLLAR__515__B[26] = __DOLLAR__procmux__DOLLAR__513__Y[26];
  assign __DOLLAR__procmux__DOLLAR__515__B[27] = __DOLLAR__procmux__DOLLAR__513__Y[27];
  assign __DOLLAR__procmux__DOLLAR__515__B[28] = __DOLLAR__procmux__DOLLAR__513__Y[28];
  assign __DOLLAR__procmux__DOLLAR__515__B[29] = __DOLLAR__procmux__DOLLAR__513__Y[29];
  assign __DOLLAR__procmux__DOLLAR__515__B[3] = __DOLLAR__procmux__DOLLAR__513__Y[3];
  assign __DOLLAR__procmux__DOLLAR__515__B[30] = __DOLLAR__procmux__DOLLAR__513__Y[30];
  assign __DOLLAR__procmux__DOLLAR__515__B[31] = __DOLLAR__procmux__DOLLAR__513__Y[31];
  assign __DOLLAR__procmux__DOLLAR__515__B[4] = __DOLLAR__procmux__DOLLAR__513__Y[4];
  assign __DOLLAR__procmux__DOLLAR__515__B[5] = __DOLLAR__procmux__DOLLAR__513__Y[5];
  assign __DOLLAR__procmux__DOLLAR__515__B[6] = __DOLLAR__procmux__DOLLAR__513__Y[6];
  assign __DOLLAR__procmux__DOLLAR__515__B[7] = __DOLLAR__procmux__DOLLAR__513__Y[7];
  assign __DOLLAR__procmux__DOLLAR__515__B[8] = __DOLLAR__procmux__DOLLAR__513__Y[8];
  assign __DOLLAR__procmux__DOLLAR__515__B[9] = __DOLLAR__procmux__DOLLAR__513__Y[9];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[0] = config_addr[24];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[1] = config_addr[25];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[2] = config_addr[26];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[3] = config_addr[27];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[4] = config_addr[28];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[5] = config_addr[29];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[6] = config_addr[30];
  assign __DOLLAR__procmux__DOLLAR__514_CMP0__A[7] = config_addr[31];
  assign __DOLLAR__procmux__DOLLAR__520__B[0] = config_data[0];
  assign __DOLLAR__procmux__DOLLAR__520__B[1] = config_data[1];
  assign __DOLLAR__procmux__DOLLAR__520__B[10] = config_data[10];
  assign __DOLLAR__procmux__DOLLAR__520__B[11] = config_data[11];
  assign __DOLLAR__procmux__DOLLAR__520__B[12] = config_data[12];
  assign __DOLLAR__procmux__DOLLAR__520__B[13] = config_data[13];
  assign __DOLLAR__procmux__DOLLAR__520__B[14] = config_data[14];
  assign __DOLLAR__procmux__DOLLAR__520__B[15] = config_data[15];
  assign __DOLLAR__procmux__DOLLAR__520__B[16] = config_data[16];
  assign __DOLLAR__procmux__DOLLAR__520__B[17] = config_data[17];
  assign __DOLLAR__procmux__DOLLAR__520__B[18] = config_data[18];
  assign __DOLLAR__procmux__DOLLAR__520__B[19] = config_data[19];
  assign __DOLLAR__procmux__DOLLAR__520__B[2] = config_data[2];
  assign __DOLLAR__procmux__DOLLAR__520__B[20] = config_data[20];
  assign __DOLLAR__procmux__DOLLAR__520__B[21] = config_data[21];
  assign __DOLLAR__procmux__DOLLAR__520__B[22] = config_data[22];
  assign __DOLLAR__procmux__DOLLAR__520__B[23] = config_data[23];
  assign __DOLLAR__procmux__DOLLAR__520__B[24] = config_data[24];
  assign __DOLLAR__procmux__DOLLAR__520__B[25] = config_data[25];
  assign __DOLLAR__procmux__DOLLAR__520__B[26] = config_data[26];
  assign __DOLLAR__procmux__DOLLAR__520__B[27] = config_data[27];
  assign __DOLLAR__procmux__DOLLAR__520__B[28] = config_data[28];
  assign __DOLLAR__procmux__DOLLAR__520__B[29] = config_data[29];
  assign __DOLLAR__procmux__DOLLAR__520__B[3] = config_data[3];
  assign __DOLLAR__procmux__DOLLAR__520__B[30] = config_data[30];
  assign __DOLLAR__procmux__DOLLAR__520__B[31] = config_data[31];
  assign __DOLLAR__procmux__DOLLAR__520__B[4] = config_data[4];
  assign __DOLLAR__procmux__DOLLAR__520__B[5] = config_data[5];
  assign __DOLLAR__procmux__DOLLAR__520__B[6] = config_data[6];
  assign __DOLLAR__procmux__DOLLAR__520__B[7] = config_data[7];
  assign __DOLLAR__procmux__DOLLAR__520__B[8] = config_data[8];
  assign __DOLLAR__procmux__DOLLAR__520__B[9] = config_data[9];
  assign __DOLLAR__procmux__DOLLAR__522__B[0] = __DOLLAR__procmux__DOLLAR__520__Y[0];
  assign __DOLLAR__procmux__DOLLAR__522__B[1] = __DOLLAR__procmux__DOLLAR__520__Y[1];
  assign __DOLLAR__procmux__DOLLAR__522__B[10] = __DOLLAR__procmux__DOLLAR__520__Y[10];
  assign __DOLLAR__procmux__DOLLAR__522__B[11] = __DOLLAR__procmux__DOLLAR__520__Y[11];
  assign __DOLLAR__procmux__DOLLAR__522__B[12] = __DOLLAR__procmux__DOLLAR__520__Y[12];
  assign __DOLLAR__procmux__DOLLAR__522__B[13] = __DOLLAR__procmux__DOLLAR__520__Y[13];
  assign __DOLLAR__procmux__DOLLAR__522__B[14] = __DOLLAR__procmux__DOLLAR__520__Y[14];
  assign __DOLLAR__procmux__DOLLAR__522__B[15] = __DOLLAR__procmux__DOLLAR__520__Y[15];
  assign __DOLLAR__procmux__DOLLAR__522__B[16] = __DOLLAR__procmux__DOLLAR__520__Y[16];
  assign __DOLLAR__procmux__DOLLAR__522__B[17] = __DOLLAR__procmux__DOLLAR__520__Y[17];
  assign __DOLLAR__procmux__DOLLAR__522__B[18] = __DOLLAR__procmux__DOLLAR__520__Y[18];
  assign __DOLLAR__procmux__DOLLAR__522__B[19] = __DOLLAR__procmux__DOLLAR__520__Y[19];
  assign __DOLLAR__procmux__DOLLAR__522__B[2] = __DOLLAR__procmux__DOLLAR__520__Y[2];
  assign __DOLLAR__procmux__DOLLAR__522__B[20] = __DOLLAR__procmux__DOLLAR__520__Y[20];
  assign __DOLLAR__procmux__DOLLAR__522__B[21] = __DOLLAR__procmux__DOLLAR__520__Y[21];
  assign __DOLLAR__procmux__DOLLAR__522__B[22] = __DOLLAR__procmux__DOLLAR__520__Y[22];
  assign __DOLLAR__procmux__DOLLAR__522__B[23] = __DOLLAR__procmux__DOLLAR__520__Y[23];
  assign __DOLLAR__procmux__DOLLAR__522__B[24] = __DOLLAR__procmux__DOLLAR__520__Y[24];
  assign __DOLLAR__procmux__DOLLAR__522__B[25] = __DOLLAR__procmux__DOLLAR__520__Y[25];
  assign __DOLLAR__procmux__DOLLAR__522__B[26] = __DOLLAR__procmux__DOLLAR__520__Y[26];
  assign __DOLLAR__procmux__DOLLAR__522__B[27] = __DOLLAR__procmux__DOLLAR__520__Y[27];
  assign __DOLLAR__procmux__DOLLAR__522__B[28] = __DOLLAR__procmux__DOLLAR__520__Y[28];
  assign __DOLLAR__procmux__DOLLAR__522__B[29] = __DOLLAR__procmux__DOLLAR__520__Y[29];
  assign __DOLLAR__procmux__DOLLAR__522__B[3] = __DOLLAR__procmux__DOLLAR__520__Y[3];
  assign __DOLLAR__procmux__DOLLAR__522__B[30] = __DOLLAR__procmux__DOLLAR__520__Y[30];
  assign __DOLLAR__procmux__DOLLAR__522__B[31] = __DOLLAR__procmux__DOLLAR__520__Y[31];
  assign __DOLLAR__procmux__DOLLAR__522__B[4] = __DOLLAR__procmux__DOLLAR__520__Y[4];
  assign __DOLLAR__procmux__DOLLAR__522__B[5] = __DOLLAR__procmux__DOLLAR__520__Y[5];
  assign __DOLLAR__procmux__DOLLAR__522__B[6] = __DOLLAR__procmux__DOLLAR__520__Y[6];
  assign __DOLLAR__procmux__DOLLAR__522__B[7] = __DOLLAR__procmux__DOLLAR__520__Y[7];
  assign __DOLLAR__procmux__DOLLAR__522__B[8] = __DOLLAR__procmux__DOLLAR__520__Y[8];
  assign __DOLLAR__procmux__DOLLAR__522__B[9] = __DOLLAR__procmux__DOLLAR__520__Y[9];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[0] = config_addr[24];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[1] = config_addr[25];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[2] = config_addr[26];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[3] = config_addr[27];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[4] = config_addr[28];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[5] = config_addr[29];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[6] = config_addr[30];
  assign __DOLLAR__procmux__DOLLAR__521_CMP0__A[7] = config_addr[31];
  assign out_0_0[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[0];
  assign out_0_0[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[1];
  assign out_0_0[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[10];
  assign out_0_0[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[11];
  assign out_0_0[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[12];
  assign out_0_0[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[13];
  assign out_0_0[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[14];
  assign out_0_0[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[15];
  assign out_0_0[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[2];
  assign out_0_0[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[3];
  assign out_0_0[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[4];
  assign out_0_0[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[5];
  assign out_0_0[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[6];
  assign out_0_0[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[7];
  assign out_0_0[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[8];
  assign out_0_0[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__238__DOLLAR__200__Y[9];
  assign out_0_1[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[0];
  assign out_0_1[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[1];
  assign out_0_1[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[10];
  assign out_0_1[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[11];
  assign out_0_1[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[12];
  assign out_0_1[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[13];
  assign out_0_1[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[14];
  assign out_0_1[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[15];
  assign out_0_1[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[2];
  assign out_0_1[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[3];
  assign out_0_1[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[4];
  assign out_0_1[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[5];
  assign out_0_1[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[6];
  assign out_0_1[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[7];
  assign out_0_1[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[8];
  assign out_0_1[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__257__DOLLAR__204__Y[9];
  assign out_0_2[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[0];
  assign out_0_2[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[1];
  assign out_0_2[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[10];
  assign out_0_2[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[11];
  assign out_0_2[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[12];
  assign out_0_2[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[13];
  assign out_0_2[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[14];
  assign out_0_2[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[15];
  assign out_0_2[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[2];
  assign out_0_2[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[3];
  assign out_0_2[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[4];
  assign out_0_2[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[5];
  assign out_0_2[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[6];
  assign out_0_2[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[7];
  assign out_0_2[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[8];
  assign out_0_2[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__276__DOLLAR__208__Y[9];
  assign out_0_3[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[0];
  assign out_0_3[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[1];
  assign out_0_3[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[10];
  assign out_0_3[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[11];
  assign out_0_3[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[12];
  assign out_0_3[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[13];
  assign out_0_3[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[14];
  assign out_0_3[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[15];
  assign out_0_3[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[2];
  assign out_0_3[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[3];
  assign out_0_3[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[4];
  assign out_0_3[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[5];
  assign out_0_3[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[6];
  assign out_0_3[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[7];
  assign out_0_3[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[8];
  assign out_0_3[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__295__DOLLAR__212__Y[9];
  assign out_0_4[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[0];
  assign out_0_4[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[1];
  assign out_0_4[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[10];
  assign out_0_4[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[11];
  assign out_0_4[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[12];
  assign out_0_4[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[13];
  assign out_0_4[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[14];
  assign out_0_4[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[15];
  assign out_0_4[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[2];
  assign out_0_4[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[3];
  assign out_0_4[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[4];
  assign out_0_4[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[5];
  assign out_0_4[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[6];
  assign out_0_4[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[7];
  assign out_0_4[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[8];
  assign out_0_4[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__314__DOLLAR__216__Y[9];
  assign out_1_0[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[0];
  assign out_1_0[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[1];
  assign out_1_0[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[10];
  assign out_1_0[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[11];
  assign out_1_0[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[12];
  assign out_1_0[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[13];
  assign out_1_0[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[14];
  assign out_1_0[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[15];
  assign out_1_0[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[2];
  assign out_1_0[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[3];
  assign out_1_0[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[4];
  assign out_1_0[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[5];
  assign out_1_0[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[6];
  assign out_1_0[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[7];
  assign out_1_0[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[8];
  assign out_1_0[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__333__DOLLAR__220__Y[9];
  assign out_1_1[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[0];
  assign out_1_1[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[1];
  assign out_1_1[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[10];
  assign out_1_1[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[11];
  assign out_1_1[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[12];
  assign out_1_1[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[13];
  assign out_1_1[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[14];
  assign out_1_1[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[15];
  assign out_1_1[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[2];
  assign out_1_1[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[3];
  assign out_1_1[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[4];
  assign out_1_1[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[5];
  assign out_1_1[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[6];
  assign out_1_1[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[7];
  assign out_1_1[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[8];
  assign out_1_1[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__352__DOLLAR__224__Y[9];
  assign out_1_2[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[0];
  assign out_1_2[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[1];
  assign out_1_2[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[10];
  assign out_1_2[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[11];
  assign out_1_2[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[12];
  assign out_1_2[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[13];
  assign out_1_2[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[14];
  assign out_1_2[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[15];
  assign out_1_2[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[2];
  assign out_1_2[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[3];
  assign out_1_2[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[4];
  assign out_1_2[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[5];
  assign out_1_2[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[6];
  assign out_1_2[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[7];
  assign out_1_2[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[8];
  assign out_1_2[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__371__DOLLAR__228__Y[9];
  assign out_1_3[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[0];
  assign out_1_3[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[1];
  assign out_1_3[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[10];
  assign out_1_3[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[11];
  assign out_1_3[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[12];
  assign out_1_3[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[13];
  assign out_1_3[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[14];
  assign out_1_3[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[15];
  assign out_1_3[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[2];
  assign out_1_3[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[3];
  assign out_1_3[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[4];
  assign out_1_3[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[5];
  assign out_1_3[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[6];
  assign out_1_3[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[7];
  assign out_1_3[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[8];
  assign out_1_3[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__390__DOLLAR__232__Y[9];
  assign out_1_4[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[0];
  assign out_1_4[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[1];
  assign out_1_4[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[10];
  assign out_1_4[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[11];
  assign out_1_4[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[12];
  assign out_1_4[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[13];
  assign out_1_4[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[14];
  assign out_1_4[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[15];
  assign out_1_4[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[2];
  assign out_1_4[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[3];
  assign out_1_4[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[4];
  assign out_1_4[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[5];
  assign out_1_4[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[6];
  assign out_1_4[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[7];
  assign out_1_4[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[8];
  assign out_1_4[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__409__DOLLAR__236__Y[9];
  assign out_2_0[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[0];
  assign out_2_0[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[1];
  assign out_2_0[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[10];
  assign out_2_0[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[11];
  assign out_2_0[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[12];
  assign out_2_0[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[13];
  assign out_2_0[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[14];
  assign out_2_0[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[15];
  assign out_2_0[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[2];
  assign out_2_0[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[3];
  assign out_2_0[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[4];
  assign out_2_0[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[5];
  assign out_2_0[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[6];
  assign out_2_0[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[7];
  assign out_2_0[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[8];
  assign out_2_0[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__428__DOLLAR__240__Y[9];
  assign out_2_1[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[0];
  assign out_2_1[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[1];
  assign out_2_1[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[10];
  assign out_2_1[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[11];
  assign out_2_1[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[12];
  assign out_2_1[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[13];
  assign out_2_1[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[14];
  assign out_2_1[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[15];
  assign out_2_1[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[2];
  assign out_2_1[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[3];
  assign out_2_1[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[4];
  assign out_2_1[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[5];
  assign out_2_1[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[6];
  assign out_2_1[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[7];
  assign out_2_1[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[8];
  assign out_2_1[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__447__DOLLAR__244__Y[9];
  assign out_2_2[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[0];
  assign out_2_2[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[1];
  assign out_2_2[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[10];
  assign out_2_2[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[11];
  assign out_2_2[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[12];
  assign out_2_2[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[13];
  assign out_2_2[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[14];
  assign out_2_2[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[15];
  assign out_2_2[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[2];
  assign out_2_2[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[3];
  assign out_2_2[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[4];
  assign out_2_2[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[5];
  assign out_2_2[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[6];
  assign out_2_2[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[7];
  assign out_2_2[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[8];
  assign out_2_2[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__466__DOLLAR__248__Y[9];
  assign out_2_3[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[0];
  assign out_2_3[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[1];
  assign out_2_3[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[10];
  assign out_2_3[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[11];
  assign out_2_3[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[12];
  assign out_2_3[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[13];
  assign out_2_3[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[14];
  assign out_2_3[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[15];
  assign out_2_3[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[2];
  assign out_2_3[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[3];
  assign out_2_3[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[4];
  assign out_2_3[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[5];
  assign out_2_3[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[6];
  assign out_2_3[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[7];
  assign out_2_3[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[8];
  assign out_2_3[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__485__DOLLAR__252__Y[9];
  assign out_2_4[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[0];
  assign out_2_4[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[1];
  assign out_2_4[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[10];
  assign out_2_4[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[11];
  assign out_2_4[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[12];
  assign out_2_4[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[13];
  assign out_2_4[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[14];
  assign out_2_4[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[15];
  assign out_2_4[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[2];
  assign out_2_4[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[3];
  assign out_2_4[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[4];
  assign out_2_4[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[5];
  assign out_2_4[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[6];
  assign out_2_4[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[7];
  assign out_2_4[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[8];
  assign out_2_4[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__504__DOLLAR__256__Y[9];
  assign out_3_0[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[0];
  assign out_3_0[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[1];
  assign out_3_0[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[10];
  assign out_3_0[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[11];
  assign out_3_0[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[12];
  assign out_3_0[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[13];
  assign out_3_0[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[14];
  assign out_3_0[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[15];
  assign out_3_0[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[2];
  assign out_3_0[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[3];
  assign out_3_0[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[4];
  assign out_3_0[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[5];
  assign out_3_0[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[6];
  assign out_3_0[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[7];
  assign out_3_0[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[8];
  assign out_3_0[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__523__DOLLAR__260__Y[9];
  assign out_3_1[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[0];
  assign out_3_1[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[1];
  assign out_3_1[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[10];
  assign out_3_1[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[11];
  assign out_3_1[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[12];
  assign out_3_1[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[13];
  assign out_3_1[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[14];
  assign out_3_1[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[15];
  assign out_3_1[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[2];
  assign out_3_1[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[3];
  assign out_3_1[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[4];
  assign out_3_1[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[5];
  assign out_3_1[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[6];
  assign out_3_1[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[7];
  assign out_3_1[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[8];
  assign out_3_1[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__542__DOLLAR__264__Y[9];
  assign out_3_2[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[0];
  assign out_3_2[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[1];
  assign out_3_2[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[10];
  assign out_3_2[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[11];
  assign out_3_2[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[12];
  assign out_3_2[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[13];
  assign out_3_2[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[14];
  assign out_3_2[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[15];
  assign out_3_2[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[2];
  assign out_3_2[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[3];
  assign out_3_2[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[4];
  assign out_3_2[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[5];
  assign out_3_2[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[6];
  assign out_3_2[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[7];
  assign out_3_2[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[8];
  assign out_3_2[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__561__DOLLAR__268__Y[9];
  assign out_3_3[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[0];
  assign out_3_3[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[1];
  assign out_3_3[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[10];
  assign out_3_3[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[11];
  assign out_3_3[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[12];
  assign out_3_3[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[13];
  assign out_3_3[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[14];
  assign out_3_3[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[15];
  assign out_3_3[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[2];
  assign out_3_3[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[3];
  assign out_3_3[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[4];
  assign out_3_3[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[5];
  assign out_3_3[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[6];
  assign out_3_3[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[7];
  assign out_3_3[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[8];
  assign out_3_3[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__580__DOLLAR__272__Y[9];
  assign out_3_4[0] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[0];
  assign out_3_4[1] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[1];
  assign out_3_4[10] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[10];
  assign out_3_4[11] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[11];
  assign out_3_4[12] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[12];
  assign out_3_4[13] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[13];
  assign out_3_4[14] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[14];
  assign out_3_4[15] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[15];
  assign out_3_4[2] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[2];
  assign out_3_4[3] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[3];
  assign out_3_4[4] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[4];
  assign out_3_4[5] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[5];
  assign out_3_4[6] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[6];
  assign out_3_4[7] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[7];
  assign out_3_4[8] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[8];
  assign out_3_4[9] = __DOLLAR__ternary__DOLLAR____DOT____FORWARD_SLASH__sb_unq1__DOT__v__COLON__599__DOLLAR__276__Y[9];

endmodule //sb_unq1

module __DOLLAR__paramod__BACKSLASH__test_shifter_unq1__BACKSLASH__DataWidth__EQUALS__16 (
  input [15:0] a,
  input [3:0] b,
  input  dir_left,
  input  is_signed,
  output [15:0] res
);
  //Wire declarations for instance '__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281' (Module shr_U21)
  wire [15:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A;
  wire [3:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B;
  wire [15:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y;
  shr_U21 __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281(
    .A(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A),
    .B(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B),
    .Y(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y)
  );

  //Wire declarations for instance '__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280' (Module sshr_U22)
  wire [15:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A;
  wire [3:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B;
  wire [15:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y;
  sshr_U22 __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280(
    .A(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A),
    .B(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B),
    .Y(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y)
  );

  //All the connections
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__S = dir_left;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__S = is_signed;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__S = dir_left;
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[0];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[1];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[10];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[11];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[12];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[13];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[14];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[15];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[2];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[3];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[4];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[5];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[6];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[7];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[8];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[9];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B[0] = b[0];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B[1] = b[1];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B[2] = b[2];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__B[3] = b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[0] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[1] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[10] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[11] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[12] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[13] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[14] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[15] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[2] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[3] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[4] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[5] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[6] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[7] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[8] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__A[9] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__281__Y[9];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[0];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[1];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[10];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[11];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[12];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[13];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[14];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[15];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[2];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[3];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[4];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[5];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[6];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[7];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[8];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__Y[9];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B[0] = b[0];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B[1] = b[1];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B[2] = b[2];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__B[3] = b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[0] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[1] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[10] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[11] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[12] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[13] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[14] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[15] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[2] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[3] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[4] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[5] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[6] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[7] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[8] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__B[9] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__280__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[0] = a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[1] = a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[10] = a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[11] = a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[12] = a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[13] = a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[14] = a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[15] = a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[2] = a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[3] = a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[4] = a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[5] = a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[6] = a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[7] = a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[8] = a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__A[9] = a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[0] = a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[1] = a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[10] = a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[11] = a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[12] = a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[13] = a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[14] = a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[15] = a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[2] = a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[3] = a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[4] = a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[5] = a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[6] = a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[7] = a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[8] = a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__279__B[9] = a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__282__Y[9];
  assign res[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[0];
  assign res[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[1];
  assign res[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[10];
  assign res[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[11];
  assign res[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[12];
  assign res[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[13];
  assign res[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[14];
  assign res[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[15];
  assign res[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[2];
  assign res[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[3];
  assign res[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[4];
  assign res[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[5];
  assign res[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[6];
  assign res[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[7];
  assign res[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[8];
  assign res[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__283__Y[9];

endmodule //__DOLLAR__paramod__BACKSLASH__test_shifter_unq1__BACKSLASH__DataWidth__EQUALS__16

module test_opt_reg (
  input  clk,
  input  clk_en,
  input [15:0] data_in,
  input  load,
  input [1:0] mode,
  output [15:0] reg_data,
  output [15:0] res,
  input  rst_n,
  input [15:0] val
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__758' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__758__ARST;
  wire  __DOLLAR__procdff__DOLLAR__758__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__758__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__758__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__758(
    .ARST(__DOLLAR__procdff__DOLLAR__758__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__758__CLK),
    .D(__DOLLAR__procdff__DOLLAR__758__D),
    .Q(__DOLLAR__procdff__DOLLAR__758__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__718' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__718__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__718__B;
  wire  __DOLLAR__procmux__DOLLAR__718__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__718__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__718(
    .A(__DOLLAR__procmux__DOLLAR__718__A),
    .B(__DOLLAR__procmux__DOLLAR__718__B),
    .S(__DOLLAR__procmux__DOLLAR__718__S),
    .Y(__DOLLAR__procmux__DOLLAR__718__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y)
  );

  //All the connections
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procdff__DOLLAR__758__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__758__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__718__S = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__S = load;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__S = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__B[0] = clk_en;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__A[0] = load;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__42__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__39__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__41__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__46__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__43__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__40__Y[0];
  assign __DOLLAR__procdff__DOLLAR__758__D[0] = __DOLLAR__procmux__DOLLAR__718__Y[0];
  assign __DOLLAR__procdff__DOLLAR__758__D[1] = __DOLLAR__procmux__DOLLAR__718__Y[1];
  assign __DOLLAR__procdff__DOLLAR__758__D[10] = __DOLLAR__procmux__DOLLAR__718__Y[10];
  assign __DOLLAR__procdff__DOLLAR__758__D[11] = __DOLLAR__procmux__DOLLAR__718__Y[11];
  assign __DOLLAR__procdff__DOLLAR__758__D[12] = __DOLLAR__procmux__DOLLAR__718__Y[12];
  assign __DOLLAR__procdff__DOLLAR__758__D[13] = __DOLLAR__procmux__DOLLAR__718__Y[13];
  assign __DOLLAR__procdff__DOLLAR__758__D[14] = __DOLLAR__procmux__DOLLAR__718__Y[14];
  assign __DOLLAR__procdff__DOLLAR__758__D[15] = __DOLLAR__procmux__DOLLAR__718__Y[15];
  assign __DOLLAR__procdff__DOLLAR__758__D[2] = __DOLLAR__procmux__DOLLAR__718__Y[2];
  assign __DOLLAR__procdff__DOLLAR__758__D[3] = __DOLLAR__procmux__DOLLAR__718__Y[3];
  assign __DOLLAR__procdff__DOLLAR__758__D[4] = __DOLLAR__procmux__DOLLAR__718__Y[4];
  assign __DOLLAR__procdff__DOLLAR__758__D[5] = __DOLLAR__procmux__DOLLAR__718__Y[5];
  assign __DOLLAR__procdff__DOLLAR__758__D[6] = __DOLLAR__procmux__DOLLAR__718__Y[6];
  assign __DOLLAR__procdff__DOLLAR__758__D[7] = __DOLLAR__procmux__DOLLAR__718__Y[7];
  assign __DOLLAR__procdff__DOLLAR__758__D[8] = __DOLLAR__procmux__DOLLAR__718__Y[8];
  assign __DOLLAR__procdff__DOLLAR__758__D[9] = __DOLLAR__procmux__DOLLAR__718__Y[9];
  assign __DOLLAR__procmux__DOLLAR__718__A[0] = __DOLLAR__procdff__DOLLAR__758__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[0] = __DOLLAR__procdff__DOLLAR__758__Q[0];
  assign reg_data[0] = __DOLLAR__procdff__DOLLAR__758__Q[0];
  assign __DOLLAR__procmux__DOLLAR__718__A[1] = __DOLLAR__procdff__DOLLAR__758__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[1] = __DOLLAR__procdff__DOLLAR__758__Q[1];
  assign reg_data[1] = __DOLLAR__procdff__DOLLAR__758__Q[1];
  assign __DOLLAR__procmux__DOLLAR__718__A[10] = __DOLLAR__procdff__DOLLAR__758__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[10] = __DOLLAR__procdff__DOLLAR__758__Q[10];
  assign reg_data[10] = __DOLLAR__procdff__DOLLAR__758__Q[10];
  assign __DOLLAR__procmux__DOLLAR__718__A[11] = __DOLLAR__procdff__DOLLAR__758__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[11] = __DOLLAR__procdff__DOLLAR__758__Q[11];
  assign reg_data[11] = __DOLLAR__procdff__DOLLAR__758__Q[11];
  assign __DOLLAR__procmux__DOLLAR__718__A[12] = __DOLLAR__procdff__DOLLAR__758__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[12] = __DOLLAR__procdff__DOLLAR__758__Q[12];
  assign reg_data[12] = __DOLLAR__procdff__DOLLAR__758__Q[12];
  assign __DOLLAR__procmux__DOLLAR__718__A[13] = __DOLLAR__procdff__DOLLAR__758__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[13] = __DOLLAR__procdff__DOLLAR__758__Q[13];
  assign reg_data[13] = __DOLLAR__procdff__DOLLAR__758__Q[13];
  assign __DOLLAR__procmux__DOLLAR__718__A[14] = __DOLLAR__procdff__DOLLAR__758__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[14] = __DOLLAR__procdff__DOLLAR__758__Q[14];
  assign reg_data[14] = __DOLLAR__procdff__DOLLAR__758__Q[14];
  assign __DOLLAR__procmux__DOLLAR__718__A[15] = __DOLLAR__procdff__DOLLAR__758__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[15] = __DOLLAR__procdff__DOLLAR__758__Q[15];
  assign reg_data[15] = __DOLLAR__procdff__DOLLAR__758__Q[15];
  assign __DOLLAR__procmux__DOLLAR__718__A[2] = __DOLLAR__procdff__DOLLAR__758__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[2] = __DOLLAR__procdff__DOLLAR__758__Q[2];
  assign reg_data[2] = __DOLLAR__procdff__DOLLAR__758__Q[2];
  assign __DOLLAR__procmux__DOLLAR__718__A[3] = __DOLLAR__procdff__DOLLAR__758__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[3] = __DOLLAR__procdff__DOLLAR__758__Q[3];
  assign reg_data[3] = __DOLLAR__procdff__DOLLAR__758__Q[3];
  assign __DOLLAR__procmux__DOLLAR__718__A[4] = __DOLLAR__procdff__DOLLAR__758__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[4] = __DOLLAR__procdff__DOLLAR__758__Q[4];
  assign reg_data[4] = __DOLLAR__procdff__DOLLAR__758__Q[4];
  assign __DOLLAR__procmux__DOLLAR__718__A[5] = __DOLLAR__procdff__DOLLAR__758__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[5] = __DOLLAR__procdff__DOLLAR__758__Q[5];
  assign reg_data[5] = __DOLLAR__procdff__DOLLAR__758__Q[5];
  assign __DOLLAR__procmux__DOLLAR__718__A[6] = __DOLLAR__procdff__DOLLAR__758__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[6] = __DOLLAR__procdff__DOLLAR__758__Q[6];
  assign reg_data[6] = __DOLLAR__procdff__DOLLAR__758__Q[6];
  assign __DOLLAR__procmux__DOLLAR__718__A[7] = __DOLLAR__procdff__DOLLAR__758__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[7] = __DOLLAR__procdff__DOLLAR__758__Q[7];
  assign reg_data[7] = __DOLLAR__procdff__DOLLAR__758__Q[7];
  assign __DOLLAR__procmux__DOLLAR__718__A[8] = __DOLLAR__procdff__DOLLAR__758__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[8] = __DOLLAR__procdff__DOLLAR__758__Q[8];
  assign reg_data[8] = __DOLLAR__procdff__DOLLAR__758__Q[8];
  assign __DOLLAR__procmux__DOLLAR__718__A[9] = __DOLLAR__procdff__DOLLAR__758__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__A[9] = __DOLLAR__procdff__DOLLAR__758__Q[9];
  assign reg_data[9] = __DOLLAR__procdff__DOLLAR__758__Q[9];
  assign __DOLLAR__procmux__DOLLAR__718__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[0];
  assign __DOLLAR__procmux__DOLLAR__718__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[1];
  assign __DOLLAR__procmux__DOLLAR__718__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[10];
  assign __DOLLAR__procmux__DOLLAR__718__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[11];
  assign __DOLLAR__procmux__DOLLAR__718__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[12];
  assign __DOLLAR__procmux__DOLLAR__718__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[13];
  assign __DOLLAR__procmux__DOLLAR__718__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[14];
  assign __DOLLAR__procmux__DOLLAR__718__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[15];
  assign __DOLLAR__procmux__DOLLAR__718__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[2];
  assign __DOLLAR__procmux__DOLLAR__718__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[3];
  assign __DOLLAR__procmux__DOLLAR__718__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[4];
  assign __DOLLAR__procmux__DOLLAR__718__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[5];
  assign __DOLLAR__procmux__DOLLAR__718__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[6];
  assign __DOLLAR__procmux__DOLLAR__718__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[7];
  assign __DOLLAR__procmux__DOLLAR__718__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[8];
  assign __DOLLAR__procmux__DOLLAR__718__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[0] = data_in[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[10] = data_in[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[11] = data_in[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[12] = data_in[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[13] = data_in[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[14] = data_in[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[15] = data_in[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[2] = data_in[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[3] = data_in[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[4] = data_in[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[5] = data_in[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[6] = data_in[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[7] = data_in[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[8] = data_in[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__A[9] = data_in[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[0] = val[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[1] = val[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[10] = val[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[11] = val[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[12] = val[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[13] = val[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[14] = val[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[15] = val[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[2] = val[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[3] = val[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[4] = val[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[5] = val[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[6] = val[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[7] = val[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[8] = val[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__38__B[9] = val[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[0] = data_in[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[10] = data_in[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[11] = data_in[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[12] = data_in[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[13] = data_in[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[14] = data_in[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[15] = data_in[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[2] = data_in[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[3] = data_in[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[4] = data_in[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[5] = data_in[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[6] = data_in[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[7] = data_in[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[8] = data_in[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__B[9] = data_in[9];
  assign res[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[0];
  assign res[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[1];
  assign res[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[10];
  assign res[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[11];
  assign res[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[12];
  assign res[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[13];
  assign res[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[14];
  assign res[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[15];
  assign res[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[2];
  assign res[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[3];
  assign res[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[4];
  assign res[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[5];
  assign res[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[6];
  assign res[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[7];
  assign res[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[8];
  assign res[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__47__Y[9];

endmodule //test_opt_reg

module test_shifter_unq1 (
  input [15:0] a,
  input [3:0] b,
  input  dir_left,
  input  is_signed,
  output [15:0] res
);
  //Wire declarations for instance '__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191' (Module shr_U21)
  wire [15:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A;
  wire [3:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B;
  wire [15:0] __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y;
  shr_U21 __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191(
    .A(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A),
    .B(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B),
    .Y(__DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y)
  );

  //Wire declarations for instance '__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190' (Module sshr_U22)
  wire [15:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A;
  wire [3:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B;
  wire [15:0] __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y;
  sshr_U22 __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190(
    .A(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A),
    .B(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B),
    .Y(__DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y)
  );

  //All the connections
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__S = dir_left;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__S = is_signed;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__S = dir_left;
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[0];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[1];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[10];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[11];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[12];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[13];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[14];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[15];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[2];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[3];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[4];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[5];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[6];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[7];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[8];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[9];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B[0] = b[0];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B[1] = b[1];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B[2] = b[2];
  assign __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__B[3] = b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[0] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[1] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[10] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[11] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[12] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[13] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[14] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[15] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[2] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[3] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[4] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[5] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[6] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[7] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[8] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__A[9] = __DOLLAR__shr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__191__Y[9];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[0];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[1];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[10];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[11];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[12];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[13];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[14];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[15];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[2];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[3];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[4];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[5];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[6];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[7];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[8];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__Y[9];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B[0] = b[0];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B[1] = b[1];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B[2] = b[2];
  assign __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__B[3] = b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[0] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[1] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[10] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[11] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[12] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[13] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[14] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[15] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[2] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[3] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[4] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[5] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[6] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[7] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[8] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__B[9] = __DOLLAR__sshr__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__190__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[0] = a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[1] = a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[10] = a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[11] = a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[12] = a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[13] = a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[14] = a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[15] = a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[2] = a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[3] = a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[4] = a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[5] = a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[6] = a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[7] = a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[8] = a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__A[9] = a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[0] = a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[1] = a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[10] = a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[11] = a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[12] = a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[13] = a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[14] = a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[15] = a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[2] = a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[3] = a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[4] = a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[5] = a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[6] = a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[7] = a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[8] = a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__70__DOLLAR__189__B[9] = a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__71__DOLLAR__192__Y[9];
  assign res[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[0];
  assign res[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[1];
  assign res[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[10];
  assign res[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[11];
  assign res[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[12];
  assign res[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[13];
  assign res[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[14];
  assign res[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[15];
  assign res[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[2];
  assign res[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[3];
  assign res[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[4];
  assign res[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[5];
  assign res[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[6];
  assign res[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[7];
  assign res[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[8];
  assign res[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_shifter_unq1__DOT__sv__COLON__85__DOLLAR__193__Y[9];

endmodule //test_shifter_unq1

module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__16 (
  input  clk,
  input  clk_en,
  input [15:0] data_in,
  input  load,
  input [1:0] mode,
  output [15:0] reg_data,
  output [15:0] res,
  input  rst_n,
  input [15:0] val
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__723' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__723__ARST;
  wire  __DOLLAR__procdff__DOLLAR__723__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__723__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__723__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__723(
    .ARST(__DOLLAR__procdff__DOLLAR__723__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__723__CLK),
    .D(__DOLLAR__procdff__DOLLAR__723__D),
    .Q(__DOLLAR__procdff__DOLLAR__723__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__356' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__356__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__356__B;
  wire  __DOLLAR__procmux__DOLLAR__356__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__356__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__356(
    .A(__DOLLAR__procmux__DOLLAR__356__A),
    .B(__DOLLAR__procmux__DOLLAR__356__B),
    .S(__DOLLAR__procmux__DOLLAR__356__S),
    .Y(__DOLLAR__procmux__DOLLAR__356__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y)
  );

  //All the connections
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procdff__DOLLAR__723__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__723__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__356__S = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__S = load;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__S = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__B[0] = clk_en;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__A[0] = load;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__349__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__346__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__348__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__353__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__350__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__347__Y[0];
  assign __DOLLAR__procdff__DOLLAR__723__D[0] = __DOLLAR__procmux__DOLLAR__356__Y[0];
  assign __DOLLAR__procdff__DOLLAR__723__D[1] = __DOLLAR__procmux__DOLLAR__356__Y[1];
  assign __DOLLAR__procdff__DOLLAR__723__D[10] = __DOLLAR__procmux__DOLLAR__356__Y[10];
  assign __DOLLAR__procdff__DOLLAR__723__D[11] = __DOLLAR__procmux__DOLLAR__356__Y[11];
  assign __DOLLAR__procdff__DOLLAR__723__D[12] = __DOLLAR__procmux__DOLLAR__356__Y[12];
  assign __DOLLAR__procdff__DOLLAR__723__D[13] = __DOLLAR__procmux__DOLLAR__356__Y[13];
  assign __DOLLAR__procdff__DOLLAR__723__D[14] = __DOLLAR__procmux__DOLLAR__356__Y[14];
  assign __DOLLAR__procdff__DOLLAR__723__D[15] = __DOLLAR__procmux__DOLLAR__356__Y[15];
  assign __DOLLAR__procdff__DOLLAR__723__D[2] = __DOLLAR__procmux__DOLLAR__356__Y[2];
  assign __DOLLAR__procdff__DOLLAR__723__D[3] = __DOLLAR__procmux__DOLLAR__356__Y[3];
  assign __DOLLAR__procdff__DOLLAR__723__D[4] = __DOLLAR__procmux__DOLLAR__356__Y[4];
  assign __DOLLAR__procdff__DOLLAR__723__D[5] = __DOLLAR__procmux__DOLLAR__356__Y[5];
  assign __DOLLAR__procdff__DOLLAR__723__D[6] = __DOLLAR__procmux__DOLLAR__356__Y[6];
  assign __DOLLAR__procdff__DOLLAR__723__D[7] = __DOLLAR__procmux__DOLLAR__356__Y[7];
  assign __DOLLAR__procdff__DOLLAR__723__D[8] = __DOLLAR__procmux__DOLLAR__356__Y[8];
  assign __DOLLAR__procdff__DOLLAR__723__D[9] = __DOLLAR__procmux__DOLLAR__356__Y[9];
  assign __DOLLAR__procmux__DOLLAR__356__A[0] = __DOLLAR__procdff__DOLLAR__723__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[0] = __DOLLAR__procdff__DOLLAR__723__Q[0];
  assign reg_data[0] = __DOLLAR__procdff__DOLLAR__723__Q[0];
  assign __DOLLAR__procmux__DOLLAR__356__A[1] = __DOLLAR__procdff__DOLLAR__723__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[1] = __DOLLAR__procdff__DOLLAR__723__Q[1];
  assign reg_data[1] = __DOLLAR__procdff__DOLLAR__723__Q[1];
  assign __DOLLAR__procmux__DOLLAR__356__A[10] = __DOLLAR__procdff__DOLLAR__723__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[10] = __DOLLAR__procdff__DOLLAR__723__Q[10];
  assign reg_data[10] = __DOLLAR__procdff__DOLLAR__723__Q[10];
  assign __DOLLAR__procmux__DOLLAR__356__A[11] = __DOLLAR__procdff__DOLLAR__723__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[11] = __DOLLAR__procdff__DOLLAR__723__Q[11];
  assign reg_data[11] = __DOLLAR__procdff__DOLLAR__723__Q[11];
  assign __DOLLAR__procmux__DOLLAR__356__A[12] = __DOLLAR__procdff__DOLLAR__723__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[12] = __DOLLAR__procdff__DOLLAR__723__Q[12];
  assign reg_data[12] = __DOLLAR__procdff__DOLLAR__723__Q[12];
  assign __DOLLAR__procmux__DOLLAR__356__A[13] = __DOLLAR__procdff__DOLLAR__723__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[13] = __DOLLAR__procdff__DOLLAR__723__Q[13];
  assign reg_data[13] = __DOLLAR__procdff__DOLLAR__723__Q[13];
  assign __DOLLAR__procmux__DOLLAR__356__A[14] = __DOLLAR__procdff__DOLLAR__723__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[14] = __DOLLAR__procdff__DOLLAR__723__Q[14];
  assign reg_data[14] = __DOLLAR__procdff__DOLLAR__723__Q[14];
  assign __DOLLAR__procmux__DOLLAR__356__A[15] = __DOLLAR__procdff__DOLLAR__723__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[15] = __DOLLAR__procdff__DOLLAR__723__Q[15];
  assign reg_data[15] = __DOLLAR__procdff__DOLLAR__723__Q[15];
  assign __DOLLAR__procmux__DOLLAR__356__A[2] = __DOLLAR__procdff__DOLLAR__723__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[2] = __DOLLAR__procdff__DOLLAR__723__Q[2];
  assign reg_data[2] = __DOLLAR__procdff__DOLLAR__723__Q[2];
  assign __DOLLAR__procmux__DOLLAR__356__A[3] = __DOLLAR__procdff__DOLLAR__723__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[3] = __DOLLAR__procdff__DOLLAR__723__Q[3];
  assign reg_data[3] = __DOLLAR__procdff__DOLLAR__723__Q[3];
  assign __DOLLAR__procmux__DOLLAR__356__A[4] = __DOLLAR__procdff__DOLLAR__723__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[4] = __DOLLAR__procdff__DOLLAR__723__Q[4];
  assign reg_data[4] = __DOLLAR__procdff__DOLLAR__723__Q[4];
  assign __DOLLAR__procmux__DOLLAR__356__A[5] = __DOLLAR__procdff__DOLLAR__723__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[5] = __DOLLAR__procdff__DOLLAR__723__Q[5];
  assign reg_data[5] = __DOLLAR__procdff__DOLLAR__723__Q[5];
  assign __DOLLAR__procmux__DOLLAR__356__A[6] = __DOLLAR__procdff__DOLLAR__723__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[6] = __DOLLAR__procdff__DOLLAR__723__Q[6];
  assign reg_data[6] = __DOLLAR__procdff__DOLLAR__723__Q[6];
  assign __DOLLAR__procmux__DOLLAR__356__A[7] = __DOLLAR__procdff__DOLLAR__723__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[7] = __DOLLAR__procdff__DOLLAR__723__Q[7];
  assign reg_data[7] = __DOLLAR__procdff__DOLLAR__723__Q[7];
  assign __DOLLAR__procmux__DOLLAR__356__A[8] = __DOLLAR__procdff__DOLLAR__723__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[8] = __DOLLAR__procdff__DOLLAR__723__Q[8];
  assign reg_data[8] = __DOLLAR__procdff__DOLLAR__723__Q[8];
  assign __DOLLAR__procmux__DOLLAR__356__A[9] = __DOLLAR__procdff__DOLLAR__723__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__A[9] = __DOLLAR__procdff__DOLLAR__723__Q[9];
  assign reg_data[9] = __DOLLAR__procdff__DOLLAR__723__Q[9];
  assign __DOLLAR__procmux__DOLLAR__356__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[0];
  assign __DOLLAR__procmux__DOLLAR__356__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[1];
  assign __DOLLAR__procmux__DOLLAR__356__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[10];
  assign __DOLLAR__procmux__DOLLAR__356__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[11];
  assign __DOLLAR__procmux__DOLLAR__356__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[12];
  assign __DOLLAR__procmux__DOLLAR__356__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[13];
  assign __DOLLAR__procmux__DOLLAR__356__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[14];
  assign __DOLLAR__procmux__DOLLAR__356__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[15];
  assign __DOLLAR__procmux__DOLLAR__356__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[2];
  assign __DOLLAR__procmux__DOLLAR__356__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[3];
  assign __DOLLAR__procmux__DOLLAR__356__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[4];
  assign __DOLLAR__procmux__DOLLAR__356__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[5];
  assign __DOLLAR__procmux__DOLLAR__356__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[6];
  assign __DOLLAR__procmux__DOLLAR__356__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[7];
  assign __DOLLAR__procmux__DOLLAR__356__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[8];
  assign __DOLLAR__procmux__DOLLAR__356__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[0] = data_in[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[10] = data_in[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[11] = data_in[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[12] = data_in[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[13] = data_in[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[14] = data_in[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[15] = data_in[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[2] = data_in[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[3] = data_in[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[4] = data_in[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[5] = data_in[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[6] = data_in[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[7] = data_in[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[8] = data_in[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__A[9] = data_in[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[0] = val[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[1] = val[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[10] = val[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[11] = val[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[12] = val[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[13] = val[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[14] = val[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[15] = val[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[2] = val[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[3] = val[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[4] = val[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[5] = val[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[6] = val[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[7] = val[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[8] = val[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__345__B[9] = val[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[0] = data_in[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[10] = data_in[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[11] = data_in[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[12] = data_in[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[13] = data_in[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[14] = data_in[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[15] = data_in[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[2] = data_in[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[3] = data_in[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[4] = data_in[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[5] = data_in[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[6] = data_in[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[7] = data_in[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[8] = data_in[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__B[9] = data_in[9];
  assign res[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[0];
  assign res[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[1];
  assign res[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[10];
  assign res[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[11];
  assign res[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[12];
  assign res[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[13];
  assign res[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[14];
  assign res[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[15];
  assign res[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[2];
  assign res[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[3];
  assign res[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[4];
  assign res[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[5];
  assign res[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[6];
  assign res[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[7];
  assign res[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[8];
  assign res[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__354__Y[9];

endmodule //__DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__16

module rtMux_U8 (
  input [0:0] A,
  input [0:0] B,
  input  S,
  output [0:0] Y
);
  //Wire declarations for instance 'mux0' (Module coreir_mux)
  wire [0:0] mux0__in0;
  wire [0:0] mux0__in1;
  wire [0:0] mux0__out;
  wire  mux0__sel;
  coreir_mux #(.width(1)) mux0(
    .in0(mux0__in0),
    .in1(mux0__in1),
    .out(mux0__out),
    .sel(mux0__sel)
  );

  //All the connections
  assign mux0__in0[0:0] = A[0:0];
  assign mux0__in1[0:0] = B[0:0];
  assign Y[0:0] = mux0__out[0:0];
  assign mux0__sel = S;

endmodule //rtMux_U8

module test_cmpr (
  input  a_msb,
  input  b_msb,
  input  diff_msb,
  input  eq,
  output  gte,
  input  is_signed,
  output  lte
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1' (Module xor_U27)
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__A;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__B;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__Y;
  xor_U27 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8' (Module xor_U27)
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__A;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__B;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__Y;
  xor_U27 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15' (Module xor_U27)
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__A;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__B;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__Y;
  xor_U27 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22' (Module xor_U27)
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__A;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__B;
  wire [0:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__Y;
  xor_U27 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__Y)
  );

  //All the connections
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__S = is_signed;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__S = is_signed;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__A[0] = a_msb;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__A[0] = a_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__A[0] = a_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__A[0] = a_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__A[0] = a_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__A[0] = a_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__A[0] = a_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__A[0] = a_msb;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__B[0] = b_msb;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__B[0] = b_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__A[0] = b_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__A[0] = b_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__B[0] = b_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__B[0] = b_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__B[0] = b_msb;
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__B[0] = b_msb;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__B[0] = diff_msb;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__B[0] = diff_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__A[0] = diff_msb;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__A[0] = diff_msb;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__B[0] = eq;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__B[0] = eq;
  assign gte = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__Y[0];
  assign lte = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__3__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__4__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__5__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__10__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__11__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__12__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__17__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__18__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__19__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__20__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__24__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__25__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__26__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__27__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__2__A[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__53__DOLLAR__1__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__9__A[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__56__DOLLAR__8__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__16__A[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__60__DOLLAR__15__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__23__A[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__63__DOLLAR__22__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__54__DOLLAR__6__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__55__DOLLAR__7__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__57__DOLLAR__13__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__66__DOLLAR__29__B[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__58__DOLLAR__14__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__61__DOLLAR__21__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__67__DOLLAR__30__B[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_cmpr__DOT__sv__COLON__64__DOLLAR__28__Y[0];

endmodule //test_cmpr

module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1 (
  input  clk,
  input  clk_en,
  input  data_in,
  input  load,
  input [1:0] mode,
  output  reg_data,
  output  res,
  input  rst_n,
  input  val
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299' (Module eq_U5)
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__A;
  wire [1:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__Y;
  eq_U5 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__728' (Module adff_U7)
  wire  __DOLLAR__procdff__DOLLAR__728__ARST;
  wire  __DOLLAR__procdff__DOLLAR__728__CLK;
  wire [0:0] __DOLLAR__procdff__DOLLAR__728__D;
  wire [0:0] __DOLLAR__procdff__DOLLAR__728__Q;
  adff_U7 #(.init(1'b0)) __DOLLAR__procdff__DOLLAR__728(
    .ARST(__DOLLAR__procdff__DOLLAR__728__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__728__CLK),
    .D(__DOLLAR__procdff__DOLLAR__728__D),
    .Q(__DOLLAR__procdff__DOLLAR__728__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__403' (Module rtMux_U8)
  wire [0:0] __DOLLAR__procmux__DOLLAR__403__A;
  wire [0:0] __DOLLAR__procmux__DOLLAR__403__B;
  wire  __DOLLAR__procmux__DOLLAR__403__S;
  wire [0:0] __DOLLAR__procmux__DOLLAR__403__Y;
  rtMux_U8 __DOLLAR__procmux__DOLLAR__403(
    .A(__DOLLAR__procmux__DOLLAR__403__A),
    .B(__DOLLAR__procmux__DOLLAR__403__B),
    .S(__DOLLAR__procmux__DOLLAR__403__S),
    .Y(__DOLLAR__procmux__DOLLAR__403__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__Y)
  );

  //All the connections
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procdff__DOLLAR__728__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__728__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__403__S = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__S = load;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__S = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__B[0] = clk_en;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__A[0] = data_in;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__B[0] = data_in;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__A[0] = load;
  assign reg_data = __DOLLAR__procdff__DOLLAR__728__Q[0];
  assign res = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__B[0] = val;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__295__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__292__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__294__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__299__A[1] = mode[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__66__DOLLAR__296__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__65__DOLLAR__293__Y[0];
  assign __DOLLAR__procdff__DOLLAR__728__D[0] = __DOLLAR__procmux__DOLLAR__403__Y[0];
  assign __DOLLAR__procmux__DOLLAR__403__A[0] = __DOLLAR__procdff__DOLLAR__728__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__76__DOLLAR__300__A[0] = __DOLLAR__procdff__DOLLAR__728__Q[0];
  assign __DOLLAR__procmux__DOLLAR__403__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg__DOT__sv__COLON__64__DOLLAR__291__Y[0];

endmodule //__DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1

module unknownBit (
  output  OUT
);
  //Wire declarations for instance 'uConst' (Module coreir_const)
  wire [0:0] uConst__out;
  coreir_const #(.value(1'bx),.width(1)) uConst(
    .out(uConst__out)
  );

  //All the connections
  assign OUT = uConst__out[0];

endmodule //unknownBit

module __DOLLAR__paramod__BACKSLASH__test_opt_reg_file__BACKSLASH__DataWidth__EQUALS__16 (
  input [7:0] cfg_a,
  input [15:0] cfg_d,
  input  cfg_en,
  input  clk,
  input  clk_en,
  input [15:0] data_in,
  input  load,
  input [2:0] mode,
  output [15:0] reg_data,
  output [15:0] res,
  input  rst_n,
  input [15:0] val
);
  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780' (Module reduce_or_U13)
  wire [1:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__Y;
  reduce_or_U13 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308' (Module eq_U18)
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__A;
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__Y;
  eq_U18 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310' (Module eq_U18)
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__A;
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__Y;
  eq_U18 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__Y)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321' (Module lt_U20)
  wire [2:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__A;
  wire [31:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B;
  wire [0:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__Y;
  lt_U20 __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321(
    .A(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__A),
    .B(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B),
    .Y(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__Y)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__724' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__724__ARST;
  wire  __DOLLAR__procdff__DOLLAR__724__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__724__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__724__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__724(
    .ARST(__DOLLAR__procdff__DOLLAR__724__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__724__CLK),
    .D(__DOLLAR__procdff__DOLLAR__724__D),
    .Q(__DOLLAR__procdff__DOLLAR__724__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__725' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__725__ARST;
  wire  __DOLLAR__procdff__DOLLAR__725__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__725__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__725__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__725(
    .ARST(__DOLLAR__procdff__DOLLAR__725__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__725__CLK),
    .D(__DOLLAR__procdff__DOLLAR__725__D),
    .Q(__DOLLAR__procdff__DOLLAR__725__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__726' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__726__ARST;
  wire  __DOLLAR__procdff__DOLLAR__726__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__726__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__726__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__726(
    .ARST(__DOLLAR__procdff__DOLLAR__726__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__726__CLK),
    .D(__DOLLAR__procdff__DOLLAR__726__D),
    .Q(__DOLLAR__procdff__DOLLAR__726__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__727' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__727__ARST;
  wire  __DOLLAR__procdff__DOLLAR__727__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__727__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__727__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__727(
    .ARST(__DOLLAR__procdff__DOLLAR__727__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__727__CLK),
    .D(__DOLLAR__procdff__DOLLAR__727__D),
    .Q(__DOLLAR__procdff__DOLLAR__727__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__359' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__359__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__359__B;
  wire  __DOLLAR__procmux__DOLLAR__359__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__359__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__359(
    .A(__DOLLAR__procmux__DOLLAR__359__A),
    .B(__DOLLAR__procmux__DOLLAR__359__B),
    .S(__DOLLAR__procmux__DOLLAR__359__S),
    .Y(__DOLLAR__procmux__DOLLAR__359__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__362' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__362__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__362__B;
  wire  __DOLLAR__procmux__DOLLAR__362__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__362__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__362(
    .A(__DOLLAR__procmux__DOLLAR__362__A),
    .B(__DOLLAR__procmux__DOLLAR__362__B),
    .S(__DOLLAR__procmux__DOLLAR__362__S),
    .Y(__DOLLAR__procmux__DOLLAR__362__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__365' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__365__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__365__B;
  wire  __DOLLAR__procmux__DOLLAR__365__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__365__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__365(
    .A(__DOLLAR__procmux__DOLLAR__365__A),
    .B(__DOLLAR__procmux__DOLLAR__365__B),
    .S(__DOLLAR__procmux__DOLLAR__365__S),
    .Y(__DOLLAR__procmux__DOLLAR__365__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__369_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__369_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__369_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__369_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__369_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__369_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__369_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__370_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__370_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__370_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__370_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__370_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__370_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__370_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__371_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__371_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__371_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__371_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__371_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__371_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__371_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__374_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__374_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__374_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__374_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__374_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__374_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__374_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__374_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__375_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__375_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__375_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__375_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__375_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__375_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__375_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__375_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__376_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__376_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__376_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__376_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__376_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__376_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__376_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__376_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__377_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__377_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__377_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__377_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__377_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__377_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__377_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__377_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__378__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__378__B;
  wire  __DOLLAR__procmux__DOLLAR__378__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__378__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__378(
    .A(__DOLLAR__procmux__DOLLAR__378__A),
    .B(__DOLLAR__procmux__DOLLAR__378__B),
    .S(__DOLLAR__procmux__DOLLAR__378__S),
    .Y(__DOLLAR__procmux__DOLLAR__378__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9(
    .OUT(__DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__379_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__379_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__379_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__379_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__379_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__379_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__379_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__379_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__382_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__382_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__382_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__382_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__382_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__382_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__382_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__382_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__383_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__383_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__383_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__383_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__383_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__383_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__383_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__383_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__391' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__391__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__391__B;
  wire  __DOLLAR__procmux__DOLLAR__391__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__391__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__391(
    .A(__DOLLAR__procmux__DOLLAR__391__A),
    .B(__DOLLAR__procmux__DOLLAR__391__B),
    .S(__DOLLAR__procmux__DOLLAR__391__S),
    .Y(__DOLLAR__procmux__DOLLAR__391__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__394' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__394__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__394__B;
  wire  __DOLLAR__procmux__DOLLAR__394__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__394__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__394(
    .A(__DOLLAR__procmux__DOLLAR__394__A),
    .B(__DOLLAR__procmux__DOLLAR__394__B),
    .S(__DOLLAR__procmux__DOLLAR__394__S),
    .Y(__DOLLAR__procmux__DOLLAR__394__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__397__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__397__B;
  wire  __DOLLAR__procmux__DOLLAR__397__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__397__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__397(
    .A(__DOLLAR__procmux__DOLLAR__397__A),
    .B(__DOLLAR__procmux__DOLLAR__397__B),
    .S(__DOLLAR__procmux__DOLLAR__397__S),
    .Y(__DOLLAR__procmux__DOLLAR__397__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9(
    .OUT(__DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__400' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__400__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__400__B;
  wire  __DOLLAR__procmux__DOLLAR__400__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__400__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__400(
    .A(__DOLLAR__procmux__DOLLAR__400__A),
    .B(__DOLLAR__procmux__DOLLAR__400__B),
    .S(__DOLLAR__procmux__DOLLAR__400__S),
    .Y(__DOLLAR__procmux__DOLLAR__400__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y)
  );

  //All the connections
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__S = __DOLLAR__procmux__DOLLAR__369_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__S = __DOLLAR__procmux__DOLLAR__371_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__S = __DOLLAR__procmux__DOLLAR__374_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__S = __DOLLAR__procmux__DOLLAR__376_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__S = __DOLLAR__procmux__DOLLAR__383_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__S = __DOLLAR__procmux__DOLLAR__382_CMP0__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[0] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[10] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[11] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[12] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[13] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[14] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[15] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[16] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[17] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[18] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[19] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[1] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[20] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[21] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[22] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[23] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[24] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[25] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[26] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[27] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[28] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[29] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[2] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[30] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[31] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[3] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[4] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[5] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[6] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[7] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[8] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__B[9] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__procdff__DOLLAR__724__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__724__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__725__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__725__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__726__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__726__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__727__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__727__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__359__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__Y[0];
  assign __DOLLAR__procmux__DOLLAR__362__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__Y[0];
  assign __DOLLAR__procmux__DOLLAR__365__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__Y[0];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__369_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__370_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__371_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__374_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__374_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__374_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__375_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__375_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__375_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__376_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__376_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__376_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__377_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__377_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__377_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__378__S = __DOLLAR__procmux__DOLLAR__379_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__378__A[0] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[10] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[11] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[12] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[13] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[14] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[15] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[1] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[2] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[3] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[4] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[5] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[6] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[7] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[8] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  assign __DOLLAR__procmux__DOLLAR__378__A[9] = __DOLLAR__procmux__DOLLAR__378__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__379_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__382_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__383_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__391__S = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__Y[0];
  assign __DOLLAR__procmux__DOLLAR__394__S = load;
  assign __DOLLAR__procmux__DOLLAR__397__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__Y[0];
  assign __DOLLAR__procmux__DOLLAR__397__B[0] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[10] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[11] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[12] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[13] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[14] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[15] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[1] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[2] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[3] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[4] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[5] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[6] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[7] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[8] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  assign __DOLLAR__procmux__DOLLAR__397__B[9] = __DOLLAR__procmux__DOLLAR__397__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  assign __DOLLAR__procmux__DOLLAR__400__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__S = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__A[0] = cfg_en;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__B[0] = clk_en;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__A[0] = load;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__328__Y[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__335__Y[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__342__Y[9];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__306__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__311__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__A[0] = __DOLLAR__procmux__DOLLAR__369_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__A[1] = __DOLLAR__procmux__DOLLAR__370_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__A[2] = __DOLLAR__procmux__DOLLAR__371_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__762__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__760__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__A[0] = __DOLLAR__procmux__DOLLAR__382_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__A[1] = __DOLLAR__procmux__DOLLAR__383_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__782__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__780__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__A[0] = __DOLLAR__procmux__DOLLAR__370_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__768__B[0] = __DOLLAR__procmux__DOLLAR__369_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__A[0] = __DOLLAR__procmux__DOLLAR__375_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__776__B[0] = __DOLLAR__procmux__DOLLAR__374_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[0] = __DOLLAR__procdff__DOLLAR__725__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[1] = __DOLLAR__procdff__DOLLAR__725__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[10] = __DOLLAR__procdff__DOLLAR__725__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[11] = __DOLLAR__procdff__DOLLAR__725__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[12] = __DOLLAR__procdff__DOLLAR__725__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[13] = __DOLLAR__procdff__DOLLAR__725__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[14] = __DOLLAR__procdff__DOLLAR__725__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[15] = __DOLLAR__procdff__DOLLAR__725__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[2] = __DOLLAR__procdff__DOLLAR__725__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[3] = __DOLLAR__procdff__DOLLAR__725__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[4] = __DOLLAR__procdff__DOLLAR__725__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[5] = __DOLLAR__procdff__DOLLAR__725__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[6] = __DOLLAR__procdff__DOLLAR__725__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[7] = __DOLLAR__procdff__DOLLAR__725__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[8] = __DOLLAR__procdff__DOLLAR__725__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__A[9] = __DOLLAR__procdff__DOLLAR__725__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[0] = __DOLLAR__procdff__DOLLAR__724__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[1] = __DOLLAR__procdff__DOLLAR__724__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[10] = __DOLLAR__procdff__DOLLAR__724__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[11] = __DOLLAR__procdff__DOLLAR__724__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[12] = __DOLLAR__procdff__DOLLAR__724__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[13] = __DOLLAR__procdff__DOLLAR__724__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[14] = __DOLLAR__procdff__DOLLAR__724__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[15] = __DOLLAR__procdff__DOLLAR__724__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[2] = __DOLLAR__procdff__DOLLAR__724__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[3] = __DOLLAR__procdff__DOLLAR__724__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[4] = __DOLLAR__procdff__DOLLAR__724__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[5] = __DOLLAR__procdff__DOLLAR__724__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[6] = __DOLLAR__procdff__DOLLAR__724__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[7] = __DOLLAR__procdff__DOLLAR__724__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[8] = __DOLLAR__procdff__DOLLAR__724__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__B[9] = __DOLLAR__procdff__DOLLAR__724__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__764__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[0] = __DOLLAR__procdff__DOLLAR__727__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[1] = __DOLLAR__procdff__DOLLAR__727__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[10] = __DOLLAR__procdff__DOLLAR__727__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[11] = __DOLLAR__procdff__DOLLAR__727__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[12] = __DOLLAR__procdff__DOLLAR__727__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[13] = __DOLLAR__procdff__DOLLAR__727__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[14] = __DOLLAR__procdff__DOLLAR__727__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[15] = __DOLLAR__procdff__DOLLAR__727__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[2] = __DOLLAR__procdff__DOLLAR__727__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[3] = __DOLLAR__procdff__DOLLAR__727__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[4] = __DOLLAR__procdff__DOLLAR__727__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[5] = __DOLLAR__procdff__DOLLAR__727__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[6] = __DOLLAR__procdff__DOLLAR__727__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[7] = __DOLLAR__procdff__DOLLAR__727__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[8] = __DOLLAR__procdff__DOLLAR__727__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__A[9] = __DOLLAR__procdff__DOLLAR__727__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[0] = __DOLLAR__procdff__DOLLAR__726__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[1] = __DOLLAR__procdff__DOLLAR__726__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[10] = __DOLLAR__procdff__DOLLAR__726__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[11] = __DOLLAR__procdff__DOLLAR__726__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[12] = __DOLLAR__procdff__DOLLAR__726__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[13] = __DOLLAR__procdff__DOLLAR__726__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[14] = __DOLLAR__procdff__DOLLAR__726__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[15] = __DOLLAR__procdff__DOLLAR__726__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[2] = __DOLLAR__procdff__DOLLAR__726__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[3] = __DOLLAR__procdff__DOLLAR__726__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[4] = __DOLLAR__procdff__DOLLAR__726__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[5] = __DOLLAR__procdff__DOLLAR__726__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[6] = __DOLLAR__procdff__DOLLAR__726__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[7] = __DOLLAR__procdff__DOLLAR__726__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[8] = __DOLLAR__procdff__DOLLAR__726__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__B[9] = __DOLLAR__procdff__DOLLAR__726__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__766__Y[9];
  assign reg_data[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[0];
  assign reg_data[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[1];
  assign reg_data[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[10];
  assign reg_data[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[11];
  assign reg_data[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[12];
  assign reg_data[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[13];
  assign reg_data[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[14];
  assign reg_data[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[15];
  assign reg_data[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[2];
  assign reg_data[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[3];
  assign reg_data[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[4];
  assign reg_data[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[5];
  assign reg_data[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[6];
  assign reg_data[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[7];
  assign reg_data[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[8];
  assign reg_data[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__770__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[0] = __DOLLAR__procdff__DOLLAR__725__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[1] = __DOLLAR__procdff__DOLLAR__725__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[10] = __DOLLAR__procdff__DOLLAR__725__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[11] = __DOLLAR__procdff__DOLLAR__725__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[12] = __DOLLAR__procdff__DOLLAR__725__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[13] = __DOLLAR__procdff__DOLLAR__725__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[14] = __DOLLAR__procdff__DOLLAR__725__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[15] = __DOLLAR__procdff__DOLLAR__725__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[2] = __DOLLAR__procdff__DOLLAR__725__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[3] = __DOLLAR__procdff__DOLLAR__725__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[4] = __DOLLAR__procdff__DOLLAR__725__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[5] = __DOLLAR__procdff__DOLLAR__725__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[6] = __DOLLAR__procdff__DOLLAR__725__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[7] = __DOLLAR__procdff__DOLLAR__725__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[8] = __DOLLAR__procdff__DOLLAR__725__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__A[9] = __DOLLAR__procdff__DOLLAR__725__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[0] = __DOLLAR__procdff__DOLLAR__724__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[1] = __DOLLAR__procdff__DOLLAR__724__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[10] = __DOLLAR__procdff__DOLLAR__724__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[11] = __DOLLAR__procdff__DOLLAR__724__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[12] = __DOLLAR__procdff__DOLLAR__724__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[13] = __DOLLAR__procdff__DOLLAR__724__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[14] = __DOLLAR__procdff__DOLLAR__724__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[15] = __DOLLAR__procdff__DOLLAR__724__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[2] = __DOLLAR__procdff__DOLLAR__724__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[3] = __DOLLAR__procdff__DOLLAR__724__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[4] = __DOLLAR__procdff__DOLLAR__724__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[5] = __DOLLAR__procdff__DOLLAR__724__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[6] = __DOLLAR__procdff__DOLLAR__724__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[7] = __DOLLAR__procdff__DOLLAR__724__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[8] = __DOLLAR__procdff__DOLLAR__724__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__B[9] = __DOLLAR__procdff__DOLLAR__724__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__772__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[0] = __DOLLAR__procdff__DOLLAR__727__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[1] = __DOLLAR__procdff__DOLLAR__727__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[10] = __DOLLAR__procdff__DOLLAR__727__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[11] = __DOLLAR__procdff__DOLLAR__727__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[12] = __DOLLAR__procdff__DOLLAR__727__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[13] = __DOLLAR__procdff__DOLLAR__727__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[14] = __DOLLAR__procdff__DOLLAR__727__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[15] = __DOLLAR__procdff__DOLLAR__727__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[2] = __DOLLAR__procdff__DOLLAR__727__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[3] = __DOLLAR__procdff__DOLLAR__727__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[4] = __DOLLAR__procdff__DOLLAR__727__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[5] = __DOLLAR__procdff__DOLLAR__727__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[6] = __DOLLAR__procdff__DOLLAR__727__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[7] = __DOLLAR__procdff__DOLLAR__727__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[8] = __DOLLAR__procdff__DOLLAR__727__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__A[9] = __DOLLAR__procdff__DOLLAR__727__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[0] = __DOLLAR__procdff__DOLLAR__726__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[1] = __DOLLAR__procdff__DOLLAR__726__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[10] = __DOLLAR__procdff__DOLLAR__726__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[11] = __DOLLAR__procdff__DOLLAR__726__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[12] = __DOLLAR__procdff__DOLLAR__726__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[13] = __DOLLAR__procdff__DOLLAR__726__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[14] = __DOLLAR__procdff__DOLLAR__726__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[15] = __DOLLAR__procdff__DOLLAR__726__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[2] = __DOLLAR__procdff__DOLLAR__726__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[3] = __DOLLAR__procdff__DOLLAR__726__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[4] = __DOLLAR__procdff__DOLLAR__726__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[5] = __DOLLAR__procdff__DOLLAR__726__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[6] = __DOLLAR__procdff__DOLLAR__726__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[7] = __DOLLAR__procdff__DOLLAR__726__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[8] = __DOLLAR__procdff__DOLLAR__726__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__B[9] = __DOLLAR__procdff__DOLLAR__726__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__774__Y[9];
  assign __DOLLAR__procmux__DOLLAR__378__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[0];
  assign __DOLLAR__procmux__DOLLAR__378__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[1];
  assign __DOLLAR__procmux__DOLLAR__378__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[10];
  assign __DOLLAR__procmux__DOLLAR__378__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[11];
  assign __DOLLAR__procmux__DOLLAR__378__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[12];
  assign __DOLLAR__procmux__DOLLAR__378__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[13];
  assign __DOLLAR__procmux__DOLLAR__378__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[14];
  assign __DOLLAR__procmux__DOLLAR__378__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[15];
  assign __DOLLAR__procmux__DOLLAR__378__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[2];
  assign __DOLLAR__procmux__DOLLAR__378__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[3];
  assign __DOLLAR__procmux__DOLLAR__378__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[4];
  assign __DOLLAR__procmux__DOLLAR__378__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[5];
  assign __DOLLAR__procmux__DOLLAR__378__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[6];
  assign __DOLLAR__procmux__DOLLAR__378__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[7];
  assign __DOLLAR__procmux__DOLLAR__378__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[8];
  assign __DOLLAR__procmux__DOLLAR__378__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__778__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[0] = __DOLLAR__procdff__DOLLAR__727__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[1] = __DOLLAR__procdff__DOLLAR__727__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[10] = __DOLLAR__procdff__DOLLAR__727__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[11] = __DOLLAR__procdff__DOLLAR__727__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[12] = __DOLLAR__procdff__DOLLAR__727__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[13] = __DOLLAR__procdff__DOLLAR__727__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[14] = __DOLLAR__procdff__DOLLAR__727__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[15] = __DOLLAR__procdff__DOLLAR__727__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[2] = __DOLLAR__procdff__DOLLAR__727__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[3] = __DOLLAR__procdff__DOLLAR__727__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[4] = __DOLLAR__procdff__DOLLAR__727__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[5] = __DOLLAR__procdff__DOLLAR__727__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[6] = __DOLLAR__procdff__DOLLAR__727__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[7] = __DOLLAR__procdff__DOLLAR__727__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[8] = __DOLLAR__procdff__DOLLAR__727__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__A[9] = __DOLLAR__procdff__DOLLAR__727__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[0] = data_in[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[1] = data_in[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[10] = data_in[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[11] = data_in[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[12] = data_in[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[13] = data_in[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[14] = data_in[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[15] = data_in[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[2] = data_in[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[3] = data_in[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[4] = data_in[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[5] = data_in[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[6] = data_in[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[7] = data_in[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[8] = data_in[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__B[9] = data_in[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__784__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__Y[9];
  assign res[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[0];
  assign res[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[1];
  assign res[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[10];
  assign res[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[11];
  assign res[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[12];
  assign res[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[13];
  assign res[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[14];
  assign res[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[15];
  assign res[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[2];
  assign res[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[3];
  assign res[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[4];
  assign res[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[5];
  assign res[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[6];
  assign res[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[7];
  assign res[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[8];
  assign res[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__786__Y[9];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__326__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__329__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__333__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__336__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__340__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__343__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__304__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__303__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__305__A[7] = cfg_a[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__A[2] = mode[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__308__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__310__A[2] = mode[2];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__330__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__327__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__337__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__334__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__344__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__341__Y[0];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__A[0] = data_in[0];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__A[1] = data_in[1];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__321__A[2] = data_in[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__307__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__312__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__309__Y[0];
  assign __DOLLAR__procdff__DOLLAR__724__D[0] = __DOLLAR__procmux__DOLLAR__359__Y[0];
  assign __DOLLAR__procdff__DOLLAR__724__D[1] = __DOLLAR__procmux__DOLLAR__359__Y[1];
  assign __DOLLAR__procdff__DOLLAR__724__D[10] = __DOLLAR__procmux__DOLLAR__359__Y[10];
  assign __DOLLAR__procdff__DOLLAR__724__D[11] = __DOLLAR__procmux__DOLLAR__359__Y[11];
  assign __DOLLAR__procdff__DOLLAR__724__D[12] = __DOLLAR__procmux__DOLLAR__359__Y[12];
  assign __DOLLAR__procdff__DOLLAR__724__D[13] = __DOLLAR__procmux__DOLLAR__359__Y[13];
  assign __DOLLAR__procdff__DOLLAR__724__D[14] = __DOLLAR__procmux__DOLLAR__359__Y[14];
  assign __DOLLAR__procdff__DOLLAR__724__D[15] = __DOLLAR__procmux__DOLLAR__359__Y[15];
  assign __DOLLAR__procdff__DOLLAR__724__D[2] = __DOLLAR__procmux__DOLLAR__359__Y[2];
  assign __DOLLAR__procdff__DOLLAR__724__D[3] = __DOLLAR__procmux__DOLLAR__359__Y[3];
  assign __DOLLAR__procdff__DOLLAR__724__D[4] = __DOLLAR__procmux__DOLLAR__359__Y[4];
  assign __DOLLAR__procdff__DOLLAR__724__D[5] = __DOLLAR__procmux__DOLLAR__359__Y[5];
  assign __DOLLAR__procdff__DOLLAR__724__D[6] = __DOLLAR__procmux__DOLLAR__359__Y[6];
  assign __DOLLAR__procdff__DOLLAR__724__D[7] = __DOLLAR__procmux__DOLLAR__359__Y[7];
  assign __DOLLAR__procdff__DOLLAR__724__D[8] = __DOLLAR__procmux__DOLLAR__359__Y[8];
  assign __DOLLAR__procdff__DOLLAR__724__D[9] = __DOLLAR__procmux__DOLLAR__359__Y[9];
  assign __DOLLAR__procmux__DOLLAR__359__A[0] = __DOLLAR__procdff__DOLLAR__724__Q[0];
  assign __DOLLAR__procmux__DOLLAR__359__A[1] = __DOLLAR__procdff__DOLLAR__724__Q[1];
  assign __DOLLAR__procmux__DOLLAR__359__A[10] = __DOLLAR__procdff__DOLLAR__724__Q[10];
  assign __DOLLAR__procmux__DOLLAR__359__A[11] = __DOLLAR__procdff__DOLLAR__724__Q[11];
  assign __DOLLAR__procmux__DOLLAR__359__A[12] = __DOLLAR__procdff__DOLLAR__724__Q[12];
  assign __DOLLAR__procmux__DOLLAR__359__A[13] = __DOLLAR__procdff__DOLLAR__724__Q[13];
  assign __DOLLAR__procmux__DOLLAR__359__A[14] = __DOLLAR__procdff__DOLLAR__724__Q[14];
  assign __DOLLAR__procmux__DOLLAR__359__A[15] = __DOLLAR__procdff__DOLLAR__724__Q[15];
  assign __DOLLAR__procmux__DOLLAR__359__A[2] = __DOLLAR__procdff__DOLLAR__724__Q[2];
  assign __DOLLAR__procmux__DOLLAR__359__A[3] = __DOLLAR__procdff__DOLLAR__724__Q[3];
  assign __DOLLAR__procmux__DOLLAR__359__A[4] = __DOLLAR__procdff__DOLLAR__724__Q[4];
  assign __DOLLAR__procmux__DOLLAR__359__A[5] = __DOLLAR__procdff__DOLLAR__724__Q[5];
  assign __DOLLAR__procmux__DOLLAR__359__A[6] = __DOLLAR__procdff__DOLLAR__724__Q[6];
  assign __DOLLAR__procmux__DOLLAR__359__A[7] = __DOLLAR__procdff__DOLLAR__724__Q[7];
  assign __DOLLAR__procmux__DOLLAR__359__A[8] = __DOLLAR__procdff__DOLLAR__724__Q[8];
  assign __DOLLAR__procmux__DOLLAR__359__A[9] = __DOLLAR__procdff__DOLLAR__724__Q[9];
  assign __DOLLAR__procdff__DOLLAR__725__D[0] = __DOLLAR__procmux__DOLLAR__362__Y[0];
  assign __DOLLAR__procdff__DOLLAR__725__D[1] = __DOLLAR__procmux__DOLLAR__362__Y[1];
  assign __DOLLAR__procdff__DOLLAR__725__D[10] = __DOLLAR__procmux__DOLLAR__362__Y[10];
  assign __DOLLAR__procdff__DOLLAR__725__D[11] = __DOLLAR__procmux__DOLLAR__362__Y[11];
  assign __DOLLAR__procdff__DOLLAR__725__D[12] = __DOLLAR__procmux__DOLLAR__362__Y[12];
  assign __DOLLAR__procdff__DOLLAR__725__D[13] = __DOLLAR__procmux__DOLLAR__362__Y[13];
  assign __DOLLAR__procdff__DOLLAR__725__D[14] = __DOLLAR__procmux__DOLLAR__362__Y[14];
  assign __DOLLAR__procdff__DOLLAR__725__D[15] = __DOLLAR__procmux__DOLLAR__362__Y[15];
  assign __DOLLAR__procdff__DOLLAR__725__D[2] = __DOLLAR__procmux__DOLLAR__362__Y[2];
  assign __DOLLAR__procdff__DOLLAR__725__D[3] = __DOLLAR__procmux__DOLLAR__362__Y[3];
  assign __DOLLAR__procdff__DOLLAR__725__D[4] = __DOLLAR__procmux__DOLLAR__362__Y[4];
  assign __DOLLAR__procdff__DOLLAR__725__D[5] = __DOLLAR__procmux__DOLLAR__362__Y[5];
  assign __DOLLAR__procdff__DOLLAR__725__D[6] = __DOLLAR__procmux__DOLLAR__362__Y[6];
  assign __DOLLAR__procdff__DOLLAR__725__D[7] = __DOLLAR__procmux__DOLLAR__362__Y[7];
  assign __DOLLAR__procdff__DOLLAR__725__D[8] = __DOLLAR__procmux__DOLLAR__362__Y[8];
  assign __DOLLAR__procdff__DOLLAR__725__D[9] = __DOLLAR__procmux__DOLLAR__362__Y[9];
  assign __DOLLAR__procmux__DOLLAR__362__A[0] = __DOLLAR__procdff__DOLLAR__725__Q[0];
  assign __DOLLAR__procmux__DOLLAR__362__A[1] = __DOLLAR__procdff__DOLLAR__725__Q[1];
  assign __DOLLAR__procmux__DOLLAR__362__A[10] = __DOLLAR__procdff__DOLLAR__725__Q[10];
  assign __DOLLAR__procmux__DOLLAR__362__A[11] = __DOLLAR__procdff__DOLLAR__725__Q[11];
  assign __DOLLAR__procmux__DOLLAR__362__A[12] = __DOLLAR__procdff__DOLLAR__725__Q[12];
  assign __DOLLAR__procmux__DOLLAR__362__A[13] = __DOLLAR__procdff__DOLLAR__725__Q[13];
  assign __DOLLAR__procmux__DOLLAR__362__A[14] = __DOLLAR__procdff__DOLLAR__725__Q[14];
  assign __DOLLAR__procmux__DOLLAR__362__A[15] = __DOLLAR__procdff__DOLLAR__725__Q[15];
  assign __DOLLAR__procmux__DOLLAR__362__A[2] = __DOLLAR__procdff__DOLLAR__725__Q[2];
  assign __DOLLAR__procmux__DOLLAR__362__A[3] = __DOLLAR__procdff__DOLLAR__725__Q[3];
  assign __DOLLAR__procmux__DOLLAR__362__A[4] = __DOLLAR__procdff__DOLLAR__725__Q[4];
  assign __DOLLAR__procmux__DOLLAR__362__A[5] = __DOLLAR__procdff__DOLLAR__725__Q[5];
  assign __DOLLAR__procmux__DOLLAR__362__A[6] = __DOLLAR__procdff__DOLLAR__725__Q[6];
  assign __DOLLAR__procmux__DOLLAR__362__A[7] = __DOLLAR__procdff__DOLLAR__725__Q[7];
  assign __DOLLAR__procmux__DOLLAR__362__A[8] = __DOLLAR__procdff__DOLLAR__725__Q[8];
  assign __DOLLAR__procmux__DOLLAR__362__A[9] = __DOLLAR__procdff__DOLLAR__725__Q[9];
  assign __DOLLAR__procdff__DOLLAR__726__D[0] = __DOLLAR__procmux__DOLLAR__365__Y[0];
  assign __DOLLAR__procdff__DOLLAR__726__D[1] = __DOLLAR__procmux__DOLLAR__365__Y[1];
  assign __DOLLAR__procdff__DOLLAR__726__D[10] = __DOLLAR__procmux__DOLLAR__365__Y[10];
  assign __DOLLAR__procdff__DOLLAR__726__D[11] = __DOLLAR__procmux__DOLLAR__365__Y[11];
  assign __DOLLAR__procdff__DOLLAR__726__D[12] = __DOLLAR__procmux__DOLLAR__365__Y[12];
  assign __DOLLAR__procdff__DOLLAR__726__D[13] = __DOLLAR__procmux__DOLLAR__365__Y[13];
  assign __DOLLAR__procdff__DOLLAR__726__D[14] = __DOLLAR__procmux__DOLLAR__365__Y[14];
  assign __DOLLAR__procdff__DOLLAR__726__D[15] = __DOLLAR__procmux__DOLLAR__365__Y[15];
  assign __DOLLAR__procdff__DOLLAR__726__D[2] = __DOLLAR__procmux__DOLLAR__365__Y[2];
  assign __DOLLAR__procdff__DOLLAR__726__D[3] = __DOLLAR__procmux__DOLLAR__365__Y[3];
  assign __DOLLAR__procdff__DOLLAR__726__D[4] = __DOLLAR__procmux__DOLLAR__365__Y[4];
  assign __DOLLAR__procdff__DOLLAR__726__D[5] = __DOLLAR__procmux__DOLLAR__365__Y[5];
  assign __DOLLAR__procdff__DOLLAR__726__D[6] = __DOLLAR__procmux__DOLLAR__365__Y[6];
  assign __DOLLAR__procdff__DOLLAR__726__D[7] = __DOLLAR__procmux__DOLLAR__365__Y[7];
  assign __DOLLAR__procdff__DOLLAR__726__D[8] = __DOLLAR__procmux__DOLLAR__365__Y[8];
  assign __DOLLAR__procdff__DOLLAR__726__D[9] = __DOLLAR__procmux__DOLLAR__365__Y[9];
  assign __DOLLAR__procmux__DOLLAR__365__A[0] = __DOLLAR__procdff__DOLLAR__726__Q[0];
  assign __DOLLAR__procmux__DOLLAR__365__A[1] = __DOLLAR__procdff__DOLLAR__726__Q[1];
  assign __DOLLAR__procmux__DOLLAR__365__A[10] = __DOLLAR__procdff__DOLLAR__726__Q[10];
  assign __DOLLAR__procmux__DOLLAR__365__A[11] = __DOLLAR__procdff__DOLLAR__726__Q[11];
  assign __DOLLAR__procmux__DOLLAR__365__A[12] = __DOLLAR__procdff__DOLLAR__726__Q[12];
  assign __DOLLAR__procmux__DOLLAR__365__A[13] = __DOLLAR__procdff__DOLLAR__726__Q[13];
  assign __DOLLAR__procmux__DOLLAR__365__A[14] = __DOLLAR__procdff__DOLLAR__726__Q[14];
  assign __DOLLAR__procmux__DOLLAR__365__A[15] = __DOLLAR__procdff__DOLLAR__726__Q[15];
  assign __DOLLAR__procmux__DOLLAR__365__A[2] = __DOLLAR__procdff__DOLLAR__726__Q[2];
  assign __DOLLAR__procmux__DOLLAR__365__A[3] = __DOLLAR__procdff__DOLLAR__726__Q[3];
  assign __DOLLAR__procmux__DOLLAR__365__A[4] = __DOLLAR__procdff__DOLLAR__726__Q[4];
  assign __DOLLAR__procmux__DOLLAR__365__A[5] = __DOLLAR__procdff__DOLLAR__726__Q[5];
  assign __DOLLAR__procmux__DOLLAR__365__A[6] = __DOLLAR__procdff__DOLLAR__726__Q[6];
  assign __DOLLAR__procmux__DOLLAR__365__A[7] = __DOLLAR__procdff__DOLLAR__726__Q[7];
  assign __DOLLAR__procmux__DOLLAR__365__A[8] = __DOLLAR__procdff__DOLLAR__726__Q[8];
  assign __DOLLAR__procmux__DOLLAR__365__A[9] = __DOLLAR__procdff__DOLLAR__726__Q[9];
  assign __DOLLAR__procdff__DOLLAR__727__D[0] = __DOLLAR__procmux__DOLLAR__391__Y[0];
  assign __DOLLAR__procdff__DOLLAR__727__D[1] = __DOLLAR__procmux__DOLLAR__391__Y[1];
  assign __DOLLAR__procdff__DOLLAR__727__D[10] = __DOLLAR__procmux__DOLLAR__391__Y[10];
  assign __DOLLAR__procdff__DOLLAR__727__D[11] = __DOLLAR__procmux__DOLLAR__391__Y[11];
  assign __DOLLAR__procdff__DOLLAR__727__D[12] = __DOLLAR__procmux__DOLLAR__391__Y[12];
  assign __DOLLAR__procdff__DOLLAR__727__D[13] = __DOLLAR__procmux__DOLLAR__391__Y[13];
  assign __DOLLAR__procdff__DOLLAR__727__D[14] = __DOLLAR__procmux__DOLLAR__391__Y[14];
  assign __DOLLAR__procdff__DOLLAR__727__D[15] = __DOLLAR__procmux__DOLLAR__391__Y[15];
  assign __DOLLAR__procdff__DOLLAR__727__D[2] = __DOLLAR__procmux__DOLLAR__391__Y[2];
  assign __DOLLAR__procdff__DOLLAR__727__D[3] = __DOLLAR__procmux__DOLLAR__391__Y[3];
  assign __DOLLAR__procdff__DOLLAR__727__D[4] = __DOLLAR__procmux__DOLLAR__391__Y[4];
  assign __DOLLAR__procdff__DOLLAR__727__D[5] = __DOLLAR__procmux__DOLLAR__391__Y[5];
  assign __DOLLAR__procdff__DOLLAR__727__D[6] = __DOLLAR__procmux__DOLLAR__391__Y[6];
  assign __DOLLAR__procdff__DOLLAR__727__D[7] = __DOLLAR__procmux__DOLLAR__391__Y[7];
  assign __DOLLAR__procdff__DOLLAR__727__D[8] = __DOLLAR__procmux__DOLLAR__391__Y[8];
  assign __DOLLAR__procdff__DOLLAR__727__D[9] = __DOLLAR__procmux__DOLLAR__391__Y[9];
  assign __DOLLAR__procmux__DOLLAR__391__A[0] = __DOLLAR__procdff__DOLLAR__727__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[0] = __DOLLAR__procdff__DOLLAR__727__Q[0];
  assign __DOLLAR__procmux__DOLLAR__391__A[1] = __DOLLAR__procdff__DOLLAR__727__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[1] = __DOLLAR__procdff__DOLLAR__727__Q[1];
  assign __DOLLAR__procmux__DOLLAR__391__A[10] = __DOLLAR__procdff__DOLLAR__727__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[10] = __DOLLAR__procdff__DOLLAR__727__Q[10];
  assign __DOLLAR__procmux__DOLLAR__391__A[11] = __DOLLAR__procdff__DOLLAR__727__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[11] = __DOLLAR__procdff__DOLLAR__727__Q[11];
  assign __DOLLAR__procmux__DOLLAR__391__A[12] = __DOLLAR__procdff__DOLLAR__727__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[12] = __DOLLAR__procdff__DOLLAR__727__Q[12];
  assign __DOLLAR__procmux__DOLLAR__391__A[13] = __DOLLAR__procdff__DOLLAR__727__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[13] = __DOLLAR__procdff__DOLLAR__727__Q[13];
  assign __DOLLAR__procmux__DOLLAR__391__A[14] = __DOLLAR__procdff__DOLLAR__727__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[14] = __DOLLAR__procdff__DOLLAR__727__Q[14];
  assign __DOLLAR__procmux__DOLLAR__391__A[15] = __DOLLAR__procdff__DOLLAR__727__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[15] = __DOLLAR__procdff__DOLLAR__727__Q[15];
  assign __DOLLAR__procmux__DOLLAR__391__A[2] = __DOLLAR__procdff__DOLLAR__727__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[2] = __DOLLAR__procdff__DOLLAR__727__Q[2];
  assign __DOLLAR__procmux__DOLLAR__391__A[3] = __DOLLAR__procdff__DOLLAR__727__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[3] = __DOLLAR__procdff__DOLLAR__727__Q[3];
  assign __DOLLAR__procmux__DOLLAR__391__A[4] = __DOLLAR__procdff__DOLLAR__727__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[4] = __DOLLAR__procdff__DOLLAR__727__Q[4];
  assign __DOLLAR__procmux__DOLLAR__391__A[5] = __DOLLAR__procdff__DOLLAR__727__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[5] = __DOLLAR__procdff__DOLLAR__727__Q[5];
  assign __DOLLAR__procmux__DOLLAR__391__A[6] = __DOLLAR__procdff__DOLLAR__727__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[6] = __DOLLAR__procdff__DOLLAR__727__Q[6];
  assign __DOLLAR__procmux__DOLLAR__391__A[7] = __DOLLAR__procdff__DOLLAR__727__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[7] = __DOLLAR__procdff__DOLLAR__727__Q[7];
  assign __DOLLAR__procmux__DOLLAR__391__A[8] = __DOLLAR__procdff__DOLLAR__727__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[8] = __DOLLAR__procdff__DOLLAR__727__Q[8];
  assign __DOLLAR__procmux__DOLLAR__391__A[9] = __DOLLAR__procdff__DOLLAR__727__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__A[9] = __DOLLAR__procdff__DOLLAR__727__Q[9];
  assign __DOLLAR__procmux__DOLLAR__359__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__359__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__359__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__359__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__359__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__359__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__359__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__359__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__359__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__359__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__359__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__359__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__359__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__359__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__359__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__359__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__362__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__362__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__362__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__362__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__362__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__362__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__362__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__362__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__362__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__362__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__362__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__362__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__362__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__362__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__362__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__362__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__365__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__365__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__365__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__365__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__365__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__365__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__365__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__365__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__365__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__365__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__365__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__365__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__365__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__365__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__365__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__365__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__369_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__370_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__371_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__374_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__374_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__375_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__375_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__376_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__376_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__377_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__377_CMP0__A[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[0] = __DOLLAR__procmux__DOLLAR__378__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[1] = __DOLLAR__procmux__DOLLAR__378__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[10] = __DOLLAR__procmux__DOLLAR__378__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[11] = __DOLLAR__procmux__DOLLAR__378__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[12] = __DOLLAR__procmux__DOLLAR__378__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[13] = __DOLLAR__procmux__DOLLAR__378__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[14] = __DOLLAR__procmux__DOLLAR__378__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[15] = __DOLLAR__procmux__DOLLAR__378__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[2] = __DOLLAR__procmux__DOLLAR__378__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[3] = __DOLLAR__procmux__DOLLAR__378__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[4] = __DOLLAR__procmux__DOLLAR__378__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[5] = __DOLLAR__procmux__DOLLAR__378__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[6] = __DOLLAR__procmux__DOLLAR__378__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[7] = __DOLLAR__procmux__DOLLAR__378__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[8] = __DOLLAR__procmux__DOLLAR__378__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__322__B[9] = __DOLLAR__procmux__DOLLAR__378__Y[9];
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__379_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__382_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__383_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__391__B[0] = __DOLLAR__procmux__DOLLAR__400__Y[0];
  assign __DOLLAR__procmux__DOLLAR__391__B[1] = __DOLLAR__procmux__DOLLAR__400__Y[1];
  assign __DOLLAR__procmux__DOLLAR__391__B[10] = __DOLLAR__procmux__DOLLAR__400__Y[10];
  assign __DOLLAR__procmux__DOLLAR__391__B[11] = __DOLLAR__procmux__DOLLAR__400__Y[11];
  assign __DOLLAR__procmux__DOLLAR__391__B[12] = __DOLLAR__procmux__DOLLAR__400__Y[12];
  assign __DOLLAR__procmux__DOLLAR__391__B[13] = __DOLLAR__procmux__DOLLAR__400__Y[13];
  assign __DOLLAR__procmux__DOLLAR__391__B[14] = __DOLLAR__procmux__DOLLAR__400__Y[14];
  assign __DOLLAR__procmux__DOLLAR__391__B[15] = __DOLLAR__procmux__DOLLAR__400__Y[15];
  assign __DOLLAR__procmux__DOLLAR__391__B[2] = __DOLLAR__procmux__DOLLAR__400__Y[2];
  assign __DOLLAR__procmux__DOLLAR__391__B[3] = __DOLLAR__procmux__DOLLAR__400__Y[3];
  assign __DOLLAR__procmux__DOLLAR__391__B[4] = __DOLLAR__procmux__DOLLAR__400__Y[4];
  assign __DOLLAR__procmux__DOLLAR__391__B[5] = __DOLLAR__procmux__DOLLAR__400__Y[5];
  assign __DOLLAR__procmux__DOLLAR__391__B[6] = __DOLLAR__procmux__DOLLAR__400__Y[6];
  assign __DOLLAR__procmux__DOLLAR__391__B[7] = __DOLLAR__procmux__DOLLAR__400__Y[7];
  assign __DOLLAR__procmux__DOLLAR__391__B[8] = __DOLLAR__procmux__DOLLAR__400__Y[8];
  assign __DOLLAR__procmux__DOLLAR__391__B[9] = __DOLLAR__procmux__DOLLAR__400__Y[9];
  assign __DOLLAR__procmux__DOLLAR__394__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__394__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__394__A[10] = data_in[10];
  assign __DOLLAR__procmux__DOLLAR__394__A[11] = data_in[11];
  assign __DOLLAR__procmux__DOLLAR__394__A[12] = data_in[12];
  assign __DOLLAR__procmux__DOLLAR__394__A[13] = data_in[13];
  assign __DOLLAR__procmux__DOLLAR__394__A[14] = data_in[14];
  assign __DOLLAR__procmux__DOLLAR__394__A[15] = data_in[15];
  assign __DOLLAR__procmux__DOLLAR__394__A[2] = data_in[2];
  assign __DOLLAR__procmux__DOLLAR__394__A[3] = data_in[3];
  assign __DOLLAR__procmux__DOLLAR__394__A[4] = data_in[4];
  assign __DOLLAR__procmux__DOLLAR__394__A[5] = data_in[5];
  assign __DOLLAR__procmux__DOLLAR__394__A[6] = data_in[6];
  assign __DOLLAR__procmux__DOLLAR__394__A[7] = data_in[7];
  assign __DOLLAR__procmux__DOLLAR__394__A[8] = data_in[8];
  assign __DOLLAR__procmux__DOLLAR__394__A[9] = data_in[9];
  assign __DOLLAR__procmux__DOLLAR__394__B[0] = val[0];
  assign __DOLLAR__procmux__DOLLAR__394__B[1] = val[1];
  assign __DOLLAR__procmux__DOLLAR__394__B[10] = val[10];
  assign __DOLLAR__procmux__DOLLAR__394__B[11] = val[11];
  assign __DOLLAR__procmux__DOLLAR__394__B[12] = val[12];
  assign __DOLLAR__procmux__DOLLAR__394__B[13] = val[13];
  assign __DOLLAR__procmux__DOLLAR__394__B[14] = val[14];
  assign __DOLLAR__procmux__DOLLAR__394__B[15] = val[15];
  assign __DOLLAR__procmux__DOLLAR__394__B[2] = val[2];
  assign __DOLLAR__procmux__DOLLAR__394__B[3] = val[3];
  assign __DOLLAR__procmux__DOLLAR__394__B[4] = val[4];
  assign __DOLLAR__procmux__DOLLAR__394__B[5] = val[5];
  assign __DOLLAR__procmux__DOLLAR__394__B[6] = val[6];
  assign __DOLLAR__procmux__DOLLAR__394__B[7] = val[7];
  assign __DOLLAR__procmux__DOLLAR__394__B[8] = val[8];
  assign __DOLLAR__procmux__DOLLAR__394__B[9] = val[9];
  assign __DOLLAR__procmux__DOLLAR__397__A[0] = __DOLLAR__procmux__DOLLAR__394__Y[0];
  assign __DOLLAR__procmux__DOLLAR__397__A[1] = __DOLLAR__procmux__DOLLAR__394__Y[1];
  assign __DOLLAR__procmux__DOLLAR__397__A[10] = __DOLLAR__procmux__DOLLAR__394__Y[10];
  assign __DOLLAR__procmux__DOLLAR__397__A[11] = __DOLLAR__procmux__DOLLAR__394__Y[11];
  assign __DOLLAR__procmux__DOLLAR__397__A[12] = __DOLLAR__procmux__DOLLAR__394__Y[12];
  assign __DOLLAR__procmux__DOLLAR__397__A[13] = __DOLLAR__procmux__DOLLAR__394__Y[13];
  assign __DOLLAR__procmux__DOLLAR__397__A[14] = __DOLLAR__procmux__DOLLAR__394__Y[14];
  assign __DOLLAR__procmux__DOLLAR__397__A[15] = __DOLLAR__procmux__DOLLAR__394__Y[15];
  assign __DOLLAR__procmux__DOLLAR__397__A[2] = __DOLLAR__procmux__DOLLAR__394__Y[2];
  assign __DOLLAR__procmux__DOLLAR__397__A[3] = __DOLLAR__procmux__DOLLAR__394__Y[3];
  assign __DOLLAR__procmux__DOLLAR__397__A[4] = __DOLLAR__procmux__DOLLAR__394__Y[4];
  assign __DOLLAR__procmux__DOLLAR__397__A[5] = __DOLLAR__procmux__DOLLAR__394__Y[5];
  assign __DOLLAR__procmux__DOLLAR__397__A[6] = __DOLLAR__procmux__DOLLAR__394__Y[6];
  assign __DOLLAR__procmux__DOLLAR__397__A[7] = __DOLLAR__procmux__DOLLAR__394__Y[7];
  assign __DOLLAR__procmux__DOLLAR__397__A[8] = __DOLLAR__procmux__DOLLAR__394__Y[8];
  assign __DOLLAR__procmux__DOLLAR__397__A[9] = __DOLLAR__procmux__DOLLAR__394__Y[9];
  assign __DOLLAR__procmux__DOLLAR__400__A[0] = __DOLLAR__procmux__DOLLAR__397__Y[0];
  assign __DOLLAR__procmux__DOLLAR__400__A[1] = __DOLLAR__procmux__DOLLAR__397__Y[1];
  assign __DOLLAR__procmux__DOLLAR__400__A[10] = __DOLLAR__procmux__DOLLAR__397__Y[10];
  assign __DOLLAR__procmux__DOLLAR__400__A[11] = __DOLLAR__procmux__DOLLAR__397__Y[11];
  assign __DOLLAR__procmux__DOLLAR__400__A[12] = __DOLLAR__procmux__DOLLAR__397__Y[12];
  assign __DOLLAR__procmux__DOLLAR__400__A[13] = __DOLLAR__procmux__DOLLAR__397__Y[13];
  assign __DOLLAR__procmux__DOLLAR__400__A[14] = __DOLLAR__procmux__DOLLAR__397__Y[14];
  assign __DOLLAR__procmux__DOLLAR__400__A[15] = __DOLLAR__procmux__DOLLAR__397__Y[15];
  assign __DOLLAR__procmux__DOLLAR__400__A[2] = __DOLLAR__procmux__DOLLAR__397__Y[2];
  assign __DOLLAR__procmux__DOLLAR__400__A[3] = __DOLLAR__procmux__DOLLAR__397__Y[3];
  assign __DOLLAR__procmux__DOLLAR__400__A[4] = __DOLLAR__procmux__DOLLAR__397__Y[4];
  assign __DOLLAR__procmux__DOLLAR__400__A[5] = __DOLLAR__procmux__DOLLAR__397__Y[5];
  assign __DOLLAR__procmux__DOLLAR__400__A[6] = __DOLLAR__procmux__DOLLAR__397__Y[6];
  assign __DOLLAR__procmux__DOLLAR__400__A[7] = __DOLLAR__procmux__DOLLAR__397__Y[7];
  assign __DOLLAR__procmux__DOLLAR__400__A[8] = __DOLLAR__procmux__DOLLAR__397__Y[8];
  assign __DOLLAR__procmux__DOLLAR__400__A[9] = __DOLLAR__procmux__DOLLAR__397__Y[9];
  assign __DOLLAR__procmux__DOLLAR__400__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__400__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__400__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__400__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__400__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__400__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__400__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__400__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__400__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__400__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__400__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__400__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__400__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__400__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__400__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__400__B[9] = cfg_d[9];

endmodule //__DOLLAR__paramod__BACKSLASH__test_opt_reg_file__BACKSLASH__DataWidth__EQUALS__16

module test_pe_comp_unq1 (
  output  carry_out,
  input [15:0] op_a,
  input [15:0] op_b,
  input [7:0] op_code,
  input  op_d_p,
  output  ovfl,
  output [15:0] res,
  output  res_p
);
  //Wire declarations for instance 'GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add' (Module __DOLLAR__paramod__BACKSLASH__test_full_add__BACKSLASH__DataWidth__EQUALS__16)
  wire [15:0] GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a;
  wire [15:0] GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b;
  wire  GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_in;
  wire  GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  wire [15:0] GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res;
  __DOLLAR__paramod__BACKSLASH__test_full_add__BACKSLASH__DataWidth__EQUALS__16 GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add(
    .a(GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a),
    .b(GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b),
    .c_in(GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_in),
    .c_out(GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out),
    .res(GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133' (Module and_U28)
  wire [15:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A;
  wire [15:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B;
  wire [15:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y;
  and_U28 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040' (Module reduce_or_U29)
  wire [4:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__Y;
  reduce_or_U29 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056' (Module reduce_or_U30)
  wire [3:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__Y;
  reduce_or_U30 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070' (Module reduce_or_U31)
  wire [14:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__Y;
  reduce_or_U31 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976' (Module reduce_or_U29)
  wire [4:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__Y;
  reduce_or_U29 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992' (Module reduce_or_U31)
  wire [14:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__Y;
  reduce_or_U31 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036' (Module reduce_or_U30)
  wire [3:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__Y;
  reduce_or_U30 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114' (Module reduce_or_U30)
  wire [3:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__Y;
  reduce_or_U30 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99' (Module eq_U32)
  wire [5:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A;
  wire [5:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__Y;
  eq_U32 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98' (Module logic_not_U33)
  wire [0:0] __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__A;
  wire [0:0] __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__Y;
  logic_not_U33 __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98(
    .A(__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__A),
    .Y(__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__Y)
  );

  //Wire declarations for instance '__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101' (Module ne_U34)
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__A;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__B;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__Y;
  ne_U34 __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101(
    .A(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__A),
    .B(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__B),
    .Y(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__Y)
  );

  //Wire declarations for instance '__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105' (Module ne_U34)
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__A;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__B;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__Y;
  ne_U34 __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105(
    .A(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__A),
    .B(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__B),
    .Y(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__Y)
  );

  //Wire declarations for instance '__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106' (Module ne_U34)
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__A;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__B;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__Y;
  ne_U34 __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106(
    .A(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__A),
    .B(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__B),
    .Y(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111' (Module not_U35)
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A;
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y;
  not_U35 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113' (Module not_U35)
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A;
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y;
  not_U35 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115' (Module not_U35)
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A;
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y;
  not_U35 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117' (Module not_U35)
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A;
  wire [15:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y;
  not_U35 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132' (Module or_U36)
  wire [15:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A;
  wire [15:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B;
  wire [15:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y;
  or_U36 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__565' (Module rtMux_U8)
  wire [0:0] __DOLLAR__procmux__DOLLAR__565__A;
  wire [0:0] __DOLLAR__procmux__DOLLAR__565__B;
  wire  __DOLLAR__procmux__DOLLAR__565__S;
  wire [0:0] __DOLLAR__procmux__DOLLAR__565__Y;
  rtMux_U8 __DOLLAR__procmux__DOLLAR__565(
    .A(__DOLLAR__procmux__DOLLAR__565__A),
    .B(__DOLLAR__procmux__DOLLAR__565__B),
    .S(__DOLLAR__procmux__DOLLAR__565__S),
    .Y(__DOLLAR__procmux__DOLLAR__565__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__567' (Module rtMux_U8)
  wire [0:0] __DOLLAR__procmux__DOLLAR__567__A;
  wire [0:0] __DOLLAR__procmux__DOLLAR__567__B;
  wire  __DOLLAR__procmux__DOLLAR__567__S;
  wire [0:0] __DOLLAR__procmux__DOLLAR__567__Y;
  rtMux_U8 __DOLLAR__procmux__DOLLAR__567(
    .A(__DOLLAR__procmux__DOLLAR__567__A),
    .B(__DOLLAR__procmux__DOLLAR__567__B),
    .S(__DOLLAR__procmux__DOLLAR__567__S),
    .Y(__DOLLAR__procmux__DOLLAR__567__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__567__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__567__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__567__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__567__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__568_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__568_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__568_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__568_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__568_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__568_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__568_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__576' (Module rtMux_U8)
  wire [0:0] __DOLLAR__procmux__DOLLAR__576__A;
  wire [0:0] __DOLLAR__procmux__DOLLAR__576__B;
  wire  __DOLLAR__procmux__DOLLAR__576__S;
  wire [0:0] __DOLLAR__procmux__DOLLAR__576__Y;
  rtMux_U8 __DOLLAR__procmux__DOLLAR__576(
    .A(__DOLLAR__procmux__DOLLAR__576__A),
    .B(__DOLLAR__procmux__DOLLAR__576__B),
    .S(__DOLLAR__procmux__DOLLAR__576__S),
    .Y(__DOLLAR__procmux__DOLLAR__576__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__578' (Module rtMux_U8)
  wire [0:0] __DOLLAR__procmux__DOLLAR__578__A;
  wire [0:0] __DOLLAR__procmux__DOLLAR__578__B;
  wire  __DOLLAR__procmux__DOLLAR__578__S;
  wire [0:0] __DOLLAR__procmux__DOLLAR__578__Y;
  rtMux_U8 __DOLLAR__procmux__DOLLAR__578(
    .A(__DOLLAR__procmux__DOLLAR__578__A),
    .B(__DOLLAR__procmux__DOLLAR__578__B),
    .S(__DOLLAR__procmux__DOLLAR__578__S),
    .Y(__DOLLAR__procmux__DOLLAR__578__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__579_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__579_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__579_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__579_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__579_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__579_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__579_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__586_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__586_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__586_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__586_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__586_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__586_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__586_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__587_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__587_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__587_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__587_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__587_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__587_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__587_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__588_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__588_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__588_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__588_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__588_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__588_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__588_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__589_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__589_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__589_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__589_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__589_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__589_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__589_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__590_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__590_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__590_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__590_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__590_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__590_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__590_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__593_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__593_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__593_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__593_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__593_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__593_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__593_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__594_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__594_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__594_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__594_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__594_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__594_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__594_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__595_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__595_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__595_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__595_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__595_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__595_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__595_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__596_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__596_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__596_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__596_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__596_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__596_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__596_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__597_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__597_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__597_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__597_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__597_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__597_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__597_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__598_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__598_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__598_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__598_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__598_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__598_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__598_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__599_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__599_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__599_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__599_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__599_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__599_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__599_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__600_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__600_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__600_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__600_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__600_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__600_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__600_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__601_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__601_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__601_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__601_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__601_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__601_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__601_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__602_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__602_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__602_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__602_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__602_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__602_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__602_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__603_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__603_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__603_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__603_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__603_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__603_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__603_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__604_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__604_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__604_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__604_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__604_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__604_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__604_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__605_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__605_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__605_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__605_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__605_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__605_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__605_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__606_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__606_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__606_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__606_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__606_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__606_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__606_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__607_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__607_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__607_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__607_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__607_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__607_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__607_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__620_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__620_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__620_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__620_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__620_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__620_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__620_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__621_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__621_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__621_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__621_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__621_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__621_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__621_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__622_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__622_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__622_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__622_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__622_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__622_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__622_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__623_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__623_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__623_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__623_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__623_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__623_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__623_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__624_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__624_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__624_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__624_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__624_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__624_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__624_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__637_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__637_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__637_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__637_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__637_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__637_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__637_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__638_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__638_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__638_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__638_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__638_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__638_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__638_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__639_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__639_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__639_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__639_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__639_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__639_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__639_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__640_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__640_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__640_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__640_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__640_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__640_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__640_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__654' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__654__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__654__B;
  wire  __DOLLAR__procmux__DOLLAR__654__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__654__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__654(
    .A(__DOLLAR__procmux__DOLLAR__654__A),
    .B(__DOLLAR__procmux__DOLLAR__654__B),
    .S(__DOLLAR__procmux__DOLLAR__654__S),
    .Y(__DOLLAR__procmux__DOLLAR__654__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__655_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__655_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__655_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__655_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__655_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__655_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__655_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__658_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__658_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__658_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__658_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__658_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__658_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__658_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__659_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__659_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__659_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__659_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__659_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__659_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__659_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__660_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__660_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__660_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__660_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__660_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__660_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__660_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__661_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__661_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__661_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__661_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__661_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__661_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__661_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__662_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__662_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__662_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__662_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__662_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__662_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__662_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__663_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__663_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__663_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__663_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__663_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__663_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__663_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__664_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__664_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__664_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__664_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__664_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__664_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__664_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__665_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__665_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__665_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__665_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__665_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__665_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__665_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__666_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__666_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__666_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__666_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__666_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__666_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__666_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__667_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__667_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__667_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__667_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__667_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__667_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__667_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__668_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__668_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__668_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__668_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__668_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__668_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__668_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__669_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__669_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__669_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__669_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__669_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__669_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__669_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__670_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__670_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__670_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__670_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__670_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__670_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__670_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__671_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__671_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__671_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__671_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__671_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__671_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__671_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0' (Module eq_U32)
  wire [5:0] __DOLLAR__procmux__DOLLAR__672_CMP0__A;
  wire [5:0] __DOLLAR__procmux__DOLLAR__672_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__672_CMP0__Y;
  eq_U32 __DOLLAR__procmux__DOLLAR__672_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__672_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__672_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__672_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97' (Module reduce_or_U37)
  wire [15:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__Y;
  reduce_or_U37 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109' (Module reduce_or_U38)
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__Y;
  reduce_or_U38 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122' (Module reduce_or_U39)
  wire [31:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__Y;
  reduce_or_U39 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125' (Module reduce_or_U37)
  wire [15:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__Y;
  reduce_or_U37 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128' (Module reduce_or_U39)
  wire [31:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__Y;
  reduce_or_U39 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131' (Module reduce_or_U40)
  wire [7:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__Y;
  reduce_or_U40 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130' (Module rtMux_U8)
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__A;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__S;
  wire [0:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__Y;
  rtMux_U8 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96' (Module xor_U41)
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A;
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B;
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y;
  xor_U41 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y)
  );

  //Wire declarations for instance '__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134' (Module xor_U41)
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A;
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B;
  wire [15:0] __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y;
  xor_U41 __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134(
    .A(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A),
    .B(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B),
    .Y(__DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y)
  );

  //Wire declarations for instance 'cmpr' (Module test_cmpr)
  wire  cmpr__a_msb;
  wire  cmpr__b_msb;
  wire  cmpr__diff_msb;
  wire  cmpr__eq;
  wire  cmpr__gte;
  wire  cmpr__is_signed;
  wire  cmpr__lte;
  test_cmpr cmpr(
    .a_msb(cmpr__a_msb),
    .b_msb(cmpr__b_msb),
    .diff_msb(cmpr__diff_msb),
    .eq(cmpr__eq),
    .gte(cmpr__gte),
    .is_signed(cmpr__is_signed),
    .lte(cmpr__lte)
  );

  //Wire declarations for instance 'test_mult_add' (Module __DOLLAR__paramod__BACKSLASH__test_mult_add__BACKSLASH__DataWidth__EQUALS__16)
  wire [15:0] test_mult_add__a;
  wire [15:0] test_mult_add__b;
  wire  test_mult_add__c_out;
  wire  test_mult_add__is_signed;
  wire [31:0] test_mult_add__res;
  __DOLLAR__paramod__BACKSLASH__test_mult_add__BACKSLASH__DataWidth__EQUALS__16 test_mult_add(
    .a(test_mult_add__a),
    .b(test_mult_add__b),
    .c_out(test_mult_add__c_out),
    .is_signed(test_mult_add__is_signed),
    .res(test_mult_add__res)
  );

  //Wire declarations for instance 'test_shifter' (Module __DOLLAR__paramod__BACKSLASH__test_shifter_unq1__BACKSLASH__DataWidth__EQUALS__16)
  wire [15:0] test_shifter__a;
  wire [3:0] test_shifter__b;
  wire  test_shifter__dir_left;
  wire  test_shifter__is_signed;
  wire [15:0] test_shifter__res;
  __DOLLAR__paramod__BACKSLASH__test_shifter_unq1__BACKSLASH__DataWidth__EQUALS__16 test_shifter(
    .a(test_shifter__a),
    .b(test_shifter__b),
    .dir_left(test_shifter__dir_left),
    .is_signed(test_shifter__is_signed),
    .res(test_shifter__res)
  );

  //All the connections
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_in = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__Y[0];
  assign carry_out = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__S = __DOLLAR__procmux__DOLLAR__597_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__S = __DOLLAR__procmux__DOLLAR__599_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__S = __DOLLAR__procmux__DOLLAR__601_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__S = __DOLLAR__procmux__DOLLAR__603_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__S = __DOLLAR__procmux__DOLLAR__605_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__S = __DOLLAR__procmux__DOLLAR__607_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__S = __DOLLAR__procmux__DOLLAR__621_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__S = __DOLLAR__procmux__DOLLAR__620_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__S = __DOLLAR__procmux__DOLLAR__624_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__S = __DOLLAR__procmux__DOLLAR__623_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__S = __DOLLAR__procmux__DOLLAR__637_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__S = __DOLLAR__procmux__DOLLAR__640_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__S = __DOLLAR__procmux__DOLLAR__639_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__S = __DOLLAR__procmux__DOLLAR__658_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__S = __DOLLAR__procmux__DOLLAR__660_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__S = __DOLLAR__procmux__DOLLAR__662_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__S = __DOLLAR__procmux__DOLLAR__664_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__S = __DOLLAR__procmux__DOLLAR__666_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__S = __DOLLAR__procmux__DOLLAR__668_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__S = __DOLLAR__procmux__DOLLAR__670_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__S = __DOLLAR__procmux__DOLLAR__672_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__S = __DOLLAR__procmux__DOLLAR__587_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__S = __DOLLAR__procmux__DOLLAR__586_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__S = __DOLLAR__procmux__DOLLAR__590_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__S = __DOLLAR__procmux__DOLLAR__589_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__S = __DOLLAR__procmux__DOLLAR__593_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__S = __DOLLAR__procmux__DOLLAR__595_CMP0__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__565__S = op_code[6];
  assign __DOLLAR__procmux__DOLLAR__567__S = __DOLLAR__procmux__DOLLAR__568_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__567__A[0] = __DOLLAR__procmux__DOLLAR__567__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__568_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__576__S = op_code[6];
  assign __DOLLAR__procmux__DOLLAR__578__S = __DOLLAR__procmux__DOLLAR__579_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__578__A[0] = __DOLLAR__procmux__DOLLAR__578__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__579_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__586_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__587_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__588_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__589_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__590_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__593_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__594_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__595_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__596_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__597_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__598_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__599_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__600_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__601_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__602_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__603_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__604_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__605_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__606_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__607_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__620_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__621_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__622_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__623_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__624_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__637_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__638_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__639_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__640_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__654__S = __DOLLAR__procmux__DOLLAR__655_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__655_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__658_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__659_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__660_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__661_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__662_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__663_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__664_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__665_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__666_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__667_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__668_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__669_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__670_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__671_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__672_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__S = op_code[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__S = op_code[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__S = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__S = cmpr__gte;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__S = cmpr__lte;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__S = op_d_p;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__S = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__S = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__Y[0];
  assign cmpr__a_msb = op_a[15];
  assign cmpr__b_msb = op_b[15];
  assign cmpr__diff_msb = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign cmpr__eq = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__A[0] = cmpr__gte;
  assign cmpr__is_signed = op_code[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__B[0] = cmpr__lte;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__A[0] = op_d_p;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__B[0] = op_d_p;
  assign ovfl = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__Y[0];
  assign res_p = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__A[0] = test_mult_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__B[0] = test_mult_add__c_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__A[0] = test_mult_add__c_out;
  assign test_mult_add__is_signed = op_code[6];
  assign test_shifter__dir_left = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__Y[0];
  assign test_shifter__is_signed = op_code[6];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[0] = __DOLLAR__procmux__DOLLAR__654__Y[0];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[1] = __DOLLAR__procmux__DOLLAR__654__Y[1];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[10] = __DOLLAR__procmux__DOLLAR__654__Y[10];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[11] = __DOLLAR__procmux__DOLLAR__654__Y[11];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[12] = __DOLLAR__procmux__DOLLAR__654__Y[12];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[13] = __DOLLAR__procmux__DOLLAR__654__Y[13];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[14] = __DOLLAR__procmux__DOLLAR__654__Y[14];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[15] = __DOLLAR__procmux__DOLLAR__654__Y[15];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[2] = __DOLLAR__procmux__DOLLAR__654__Y[2];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[3] = __DOLLAR__procmux__DOLLAR__654__Y[3];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[4] = __DOLLAR__procmux__DOLLAR__654__Y[4];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[5] = __DOLLAR__procmux__DOLLAR__654__Y[5];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[6] = __DOLLAR__procmux__DOLLAR__654__Y[6];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[7] = __DOLLAR__procmux__DOLLAR__654__Y[7];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[8] = __DOLLAR__procmux__DOLLAR__654__Y[8];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__a[9] = __DOLLAR__procmux__DOLLAR__654__Y[9];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[0];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[1];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[10];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[11];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[12];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[13];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[14];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[15];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[2];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[3];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[4];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[5];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[6];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[7];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[8];
  assign GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__b[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[1] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[1] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[1] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[10] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[10] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[10] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[11] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[11] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[11] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[12] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[12] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[12] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[13] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[13] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[13] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[14] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[14] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[14] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[15] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[15] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__A[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__B[0] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[15] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[2] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[2] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[2] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[3] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[3] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[3] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[4] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[4] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[4] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[5] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[5] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[5] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[6] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[6] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[6] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[7] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[7] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[7] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[8] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[8] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[8] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__A[9] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__B[9] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__A[9] = GEN_ADD__LEFT_BRACKET__0__RIGHT_BRACKET____DOT__full_add__res[9];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__B[0] = __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__Y[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__102__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__A[0] = __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__B[0] = __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__107__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__B[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__123__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__B[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__129__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[0] = op_a[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[1] = op_a[1];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[10] = op_a[10];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[11] = op_a[11];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[12] = op_a[12];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[13] = op_a[13];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[14] = op_a[14];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[15] = op_a[15];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[2] = op_a[2];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[3] = op_a[3];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[4] = op_a[4];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[5] = op_a[5];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[6] = op_a[6];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[7] = op_a[7];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[8] = op_a[8];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__A[9] = op_a[9];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[0] = op_b[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[1] = op_b[1];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[10] = op_b[10];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[11] = op_b[11];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[12] = op_b[12];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[13] = op_b[13];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[14] = op_b[14];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[15] = op_b[15];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[2] = op_b[2];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[3] = op_b[3];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[4] = op_b[4];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[5] = op_b[5];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[6] = op_b[6];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[7] = op_b[7];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[8] = op_b[8];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__B[9] = op_b[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[1] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[10] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[11] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[12] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[13] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[14] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[15] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[2] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[3] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[4] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[5] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[6] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[7] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[8] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__A[9] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__344__DOLLAR__133__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A[0] = __DOLLAR__procmux__DOLLAR__620_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A[1] = __DOLLAR__procmux__DOLLAR__621_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A[2] = __DOLLAR__procmux__DOLLAR__622_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A[3] = __DOLLAR__procmux__DOLLAR__623_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__A[4] = __DOLLAR__procmux__DOLLAR__624_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1042__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1040__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A[0] = __DOLLAR__procmux__DOLLAR__637_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A[1] = __DOLLAR__procmux__DOLLAR__638_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A[2] = __DOLLAR__procmux__DOLLAR__639_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__A[3] = __DOLLAR__procmux__DOLLAR__640_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1058__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1056__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[0] = __DOLLAR__procmux__DOLLAR__658_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[1] = __DOLLAR__procmux__DOLLAR__659_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[10] = __DOLLAR__procmux__DOLLAR__668_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[11] = __DOLLAR__procmux__DOLLAR__669_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[12] = __DOLLAR__procmux__DOLLAR__670_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[13] = __DOLLAR__procmux__DOLLAR__671_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[14] = __DOLLAR__procmux__DOLLAR__672_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[2] = __DOLLAR__procmux__DOLLAR__660_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[3] = __DOLLAR__procmux__DOLLAR__661_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[4] = __DOLLAR__procmux__DOLLAR__662_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[5] = __DOLLAR__procmux__DOLLAR__663_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[6] = __DOLLAR__procmux__DOLLAR__664_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[7] = __DOLLAR__procmux__DOLLAR__665_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[8] = __DOLLAR__procmux__DOLLAR__666_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__A[9] = __DOLLAR__procmux__DOLLAR__667_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1072__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1070__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A[0] = __DOLLAR__procmux__DOLLAR__586_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A[1] = __DOLLAR__procmux__DOLLAR__587_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A[2] = __DOLLAR__procmux__DOLLAR__588_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A[3] = __DOLLAR__procmux__DOLLAR__589_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__A[4] = __DOLLAR__procmux__DOLLAR__590_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__978__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__976__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[0] = __DOLLAR__procmux__DOLLAR__593_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[1] = __DOLLAR__procmux__DOLLAR__594_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[10] = __DOLLAR__procmux__DOLLAR__603_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[11] = __DOLLAR__procmux__DOLLAR__604_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[12] = __DOLLAR__procmux__DOLLAR__605_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[13] = __DOLLAR__procmux__DOLLAR__606_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[14] = __DOLLAR__procmux__DOLLAR__607_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[2] = __DOLLAR__procmux__DOLLAR__595_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[3] = __DOLLAR__procmux__DOLLAR__596_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[4] = __DOLLAR__procmux__DOLLAR__597_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[5] = __DOLLAR__procmux__DOLLAR__598_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[6] = __DOLLAR__procmux__DOLLAR__599_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[7] = __DOLLAR__procmux__DOLLAR__600_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[8] = __DOLLAR__procmux__DOLLAR__601_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__A[9] = __DOLLAR__procmux__DOLLAR__602_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__994__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__992__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__A[0] = __DOLLAR__procmux__DOLLAR__594_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__B[0] = __DOLLAR__procmux__DOLLAR__593_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1000__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__A[0] = __DOLLAR__procmux__DOLLAR__598_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__B[0] = __DOLLAR__procmux__DOLLAR__597_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1008__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__A[0] = __DOLLAR__procmux__DOLLAR__602_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__B[0] = __DOLLAR__procmux__DOLLAR__601_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1020__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__A[0] = __DOLLAR__procmux__DOLLAR__606_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1028__B[0] = __DOLLAR__procmux__DOLLAR__605_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__A[0] = __DOLLAR__procmux__DOLLAR__638_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1066__B[0] = __DOLLAR__procmux__DOLLAR__637_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__A[0] = __DOLLAR__procmux__DOLLAR__659_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__B[0] = __DOLLAR__procmux__DOLLAR__658_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1078__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__A[0] = __DOLLAR__procmux__DOLLAR__663_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__B[0] = __DOLLAR__procmux__DOLLAR__662_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1086__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__A[0] = __DOLLAR__procmux__DOLLAR__667_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__B[0] = __DOLLAR__procmux__DOLLAR__666_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1098__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__A[0] = __DOLLAR__procmux__DOLLAR__671_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1106__B[0] = __DOLLAR__procmux__DOLLAR__670_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__A[0] = __DOLLAR__procmux__DOLLAR__596_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__A[1] = __DOLLAR__procmux__DOLLAR__595_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1012__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__A[0] = __DOLLAR__procmux__DOLLAR__604_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1032__A[1] = __DOLLAR__procmux__DOLLAR__603_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A[0] = __DOLLAR__procmux__DOLLAR__600_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1036__A[1] = __DOLLAR__procmux__DOLLAR__599_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__A[0] = __DOLLAR__procmux__DOLLAR__622_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__A[1] = __DOLLAR__procmux__DOLLAR__621_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1052__A[2] = __DOLLAR__procmux__DOLLAR__620_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__A[0] = __DOLLAR__procmux__DOLLAR__661_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__A[1] = __DOLLAR__procmux__DOLLAR__660_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1090__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__A[0] = __DOLLAR__procmux__DOLLAR__669_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1110__A[1] = __DOLLAR__procmux__DOLLAR__668_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A[0] = __DOLLAR__procmux__DOLLAR__665_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1114__A[1] = __DOLLAR__procmux__DOLLAR__664_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__A[0] = __DOLLAR__procmux__DOLLAR__588_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__A[1] = __DOLLAR__procmux__DOLLAR__587_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__988__A[2] = __DOLLAR__procmux__DOLLAR__586_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__998__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__996__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1002__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1004__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1006__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1010__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1014__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1016__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1018__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1022__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__B[0] = op_a[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1024__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1026__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1030__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1038__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1034__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1044__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1046__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1048__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1054__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1050__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[1] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[10] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[11] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[12] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[13] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[14] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[15] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[2] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[3] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[4] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[5] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[6] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[7] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[8] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__A[9] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[1] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[10] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[11] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[12] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[13] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[14] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[15] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[2] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[3] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[4] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[5] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[6] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[7] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[8] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__B[9] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1060__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[0] = op_b[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[1] = op_b[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[10] = op_b[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[11] = op_b[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[12] = op_b[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[13] = op_b[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[14] = op_b[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[15] = op_b[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[2] = op_b[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[3] = op_b[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[4] = op_b[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[5] = op_b[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[6] = op_b[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[7] = op_b[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[8] = op_b[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__A[9] = op_b[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[1] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[10] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[11] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[12] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[13] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[14] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[15] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[2] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[3] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[4] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[5] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[6] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[7] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[8] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__B[9] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1062__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1068__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1064__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[1] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[10] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[11] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[12] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[13] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[14] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[15] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[2] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[3] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[4] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[5] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[6] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[7] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[8] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__B[9] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1074__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[0] = test_mult_add__res[16];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[1] = test_mult_add__res[17];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[10] = test_mult_add__res[26];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[11] = test_mult_add__res[27];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[12] = test_mult_add__res[28];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[13] = test_mult_add__res[29];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[14] = test_mult_add__res[30];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[15] = test_mult_add__res[31];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[2] = test_mult_add__res[18];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[3] = test_mult_add__res[19];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[4] = test_mult_add__res[20];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[5] = test_mult_add__res[21];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[6] = test_mult_add__res[22];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[7] = test_mult_add__res[23];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[8] = test_mult_add__res[24];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__A[9] = test_mult_add__res[25];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[1] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[10] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[11] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[12] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[13] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[14] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[15] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[2] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[3] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[4] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[5] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[6] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[7] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[8] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__B[9] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1076__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1080__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[0] = test_mult_add__res[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[1] = test_mult_add__res[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[10] = test_mult_add__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[11] = test_mult_add__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[12] = test_mult_add__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[13] = test_mult_add__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[14] = test_mult_add__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[15] = test_mult_add__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[2] = test_mult_add__res[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[3] = test_mult_add__res[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[4] = test_mult_add__res[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[5] = test_mult_add__res[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[6] = test_mult_add__res[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[7] = test_mult_add__res[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[8] = test_mult_add__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__A[9] = test_mult_add__res[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[0] = test_mult_add__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[1] = test_mult_add__res[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[10] = test_mult_add__res[18];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[11] = test_mult_add__res[19];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[12] = test_mult_add__res[20];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[13] = test_mult_add__res[21];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[14] = test_mult_add__res[22];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[15] = test_mult_add__res[23];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[2] = test_mult_add__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[3] = test_mult_add__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[4] = test_mult_add__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[5] = test_mult_add__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[6] = test_mult_add__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[7] = test_mult_add__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[8] = test_mult_add__res[16];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__B[9] = test_mult_add__res[17];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1082__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[0] = test_shifter__res[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[1] = test_shifter__res[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[10] = test_shifter__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[11] = test_shifter__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[12] = test_shifter__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[13] = test_shifter__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[14] = test_shifter__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[15] = test_shifter__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[2] = test_shifter__res[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[3] = test_shifter__res[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[4] = test_shifter__res[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[5] = test_shifter__res[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[6] = test_shifter__res[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[7] = test_shifter__res[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[8] = test_shifter__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__A[9] = test_shifter__res[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[0] = test_shifter__res[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[1] = test_shifter__res[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[10] = test_shifter__res[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[11] = test_shifter__res[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[12] = test_shifter__res[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[13] = test_shifter__res[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[14] = test_shifter__res[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[15] = test_shifter__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[2] = test_shifter__res[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[3] = test_shifter__res[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[4] = test_shifter__res[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[5] = test_shifter__res[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[6] = test_shifter__res[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[7] = test_shifter__res[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[8] = test_shifter__res[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__B[9] = test_shifter__res[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1084__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1088__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1092__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[0] = op_b[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[1] = op_b[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[10] = op_b[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[11] = op_b[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[12] = op_b[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[13] = op_b[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[14] = op_b[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[15] = op_b[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[2] = op_b[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[3] = op_b[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[4] = op_b[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[5] = op_b[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[6] = op_b[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[7] = op_b[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[8] = op_b[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__A[9] = op_b[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1094__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1096__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1100__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1102__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[0] = op_a[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[1] = op_a[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[10] = op_a[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[11] = op_a[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[12] = op_a[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[13] = op_a[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[14] = op_a[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[15] = op_a[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[2] = op_a[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[3] = op_a[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[4] = op_a[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[5] = op_a[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[6] = op_a[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[7] = op_a[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[8] = op_a[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__A[9] = op_a[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1104__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1108__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1112__Y[9];
  assign res[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[0];
  assign res[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[1];
  assign res[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[10];
  assign res[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[11];
  assign res[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[12];
  assign res[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[13];
  assign res[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[14];
  assign res[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[15];
  assign res[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[2];
  assign res[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[3];
  assign res[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[4];
  assign res[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[5];
  assign res[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[6];
  assign res[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[7];
  assign res[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[8];
  assign res[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1116__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__B[0] = __DOLLAR__procmux__DOLLAR__578__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__980__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__B[0] = __DOLLAR__procmux__DOLLAR__567__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__982__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__984__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__273__DOLLAR__112__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__990__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__986__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[0] = op_code[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[1] = op_code[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[2] = op_code[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[3] = op_code[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[4] = op_code[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__223__DOLLAR__99__A[5] = op_code[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__A[0] = op_a[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__243__DOLLAR__100__B[0] = op_b[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__A[0] = op_a[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__315__DOLLAR__120__B[0] = op_b[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__A[0] = op_a[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__326__DOLLAR__126__B[0] = op_b[15];
  assign __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__98__A[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__Y[0];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__244__DOLLAR__101__A[0] = op_a[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__A[0] = op_a[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__105__B[0] = op_b[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__248__DOLLAR__106__A[0] = op_a[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[0] = op_b[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[1] = op_b[1];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[10] = op_b[10];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[11] = op_b[11];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[12] = op_b[12];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[13] = op_b[13];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[14] = op_b[14];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[15] = op_b[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[2] = op_b[2];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[3] = op_b[3];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[4] = op_b[4];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[5] = op_b[5];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[6] = op_b[6];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[7] = op_b[7];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[8] = op_b[8];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__271__DOLLAR__111__A[9] = op_b[9];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[0] = op_a[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[1] = op_a[1];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[10] = op_a[10];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[11] = op_a[11];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[12] = op_a[12];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[13] = op_a[13];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[14] = op_a[14];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[15] = op_a[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[2] = op_a[2];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[3] = op_a[3];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[4] = op_a[4];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[5] = op_a[5];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[6] = op_a[6];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[7] = op_a[7];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[8] = op_a[8];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__A[9] = op_a[9];
  assign __DOLLAR__procmux__DOLLAR__654__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[0];
  assign __DOLLAR__procmux__DOLLAR__654__B[1] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[1];
  assign __DOLLAR__procmux__DOLLAR__654__B[10] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[10];
  assign __DOLLAR__procmux__DOLLAR__654__B[11] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[11];
  assign __DOLLAR__procmux__DOLLAR__654__B[12] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[12];
  assign __DOLLAR__procmux__DOLLAR__654__B[13] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[13];
  assign __DOLLAR__procmux__DOLLAR__654__B[14] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[14];
  assign __DOLLAR__procmux__DOLLAR__654__B[15] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[15];
  assign __DOLLAR__procmux__DOLLAR__654__B[2] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[2];
  assign __DOLLAR__procmux__DOLLAR__654__B[3] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[3];
  assign __DOLLAR__procmux__DOLLAR__654__B[4] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[4];
  assign __DOLLAR__procmux__DOLLAR__654__B[5] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[5];
  assign __DOLLAR__procmux__DOLLAR__654__B[6] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[6];
  assign __DOLLAR__procmux__DOLLAR__654__B[7] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[7];
  assign __DOLLAR__procmux__DOLLAR__654__B[8] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[8];
  assign __DOLLAR__procmux__DOLLAR__654__B[9] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__276__DOLLAR__113__Y[9];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[0] = op_b[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[1] = op_b[1];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[10] = op_b[10];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[11] = op_b[11];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[12] = op_b[12];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[13] = op_b[13];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[14] = op_b[14];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[15] = op_b[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[2] = op_b[2];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[3] = op_b[3];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[4] = op_b[4];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[5] = op_b[5];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[6] = op_b[6];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[7] = op_b[7];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[8] = op_b[8];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__287__DOLLAR__115__A[9] = op_b[9];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[0] = op_b[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[1] = op_b[1];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[10] = op_b[10];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[11] = op_b[11];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[12] = op_b[12];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[13] = op_b[13];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[14] = op_b[14];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[15] = op_b[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[2] = op_b[2];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[3] = op_b[3];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[4] = op_b[4];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[5] = op_b[5];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[6] = op_b[6];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[7] = op_b[7];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[8] = op_b[8];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__293__DOLLAR__117__A[9] = op_b[9];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__121__A[0] = test_mult_add__res[15];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__127__A[0] = test_mult_add__res[15];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[0] = op_a[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[1] = op_a[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[10] = op_a[10];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[11] = op_a[11];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[12] = op_a[12];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[13] = op_a[13];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[14] = op_a[14];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[15] = op_a[15];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[2] = op_a[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[3] = op_a[3];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[4] = op_a[4];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[5] = op_a[5];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[6] = op_a[6];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[7] = op_a[7];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[8] = op_a[8];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__A[9] = op_a[9];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[0] = op_b[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[1] = op_b[1];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[10] = op_b[10];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[11] = op_b[11];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[12] = op_b[12];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[13] = op_b[13];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[14] = op_b[14];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[15] = op_b[15];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[2] = op_b[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[3] = op_b[3];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[4] = op_b[4];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[5] = op_b[5];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[6] = op_b[6];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[7] = op_b[7];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[8] = op_b[8];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__341__DOLLAR__132__B[9] = op_b[9];
  assign __DOLLAR__procmux__DOLLAR__565__A[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__Y[0];
  assign __DOLLAR__procmux__DOLLAR__565__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__Y[0];
  assign __DOLLAR__procmux__DOLLAR__567__B[0] = __DOLLAR__procmux__DOLLAR__565__Y[0];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__568_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__576__A[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__Y[0];
  assign __DOLLAR__procmux__DOLLAR__576__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__Y[0];
  assign __DOLLAR__procmux__DOLLAR__578__B[0] = __DOLLAR__procmux__DOLLAR__576__Y[0];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__579_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__586_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__587_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__588_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__589_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__590_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__593_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__594_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__595_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__596_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__597_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__598_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__599_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__600_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__601_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__602_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__603_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__604_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__605_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__606_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__607_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__620_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__621_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__622_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__623_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__624_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__637_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__638_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__639_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__640_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__654__A[0] = op_a[0];
  assign __DOLLAR__procmux__DOLLAR__654__A[1] = op_a[1];
  assign __DOLLAR__procmux__DOLLAR__654__A[10] = op_a[10];
  assign __DOLLAR__procmux__DOLLAR__654__A[11] = op_a[11];
  assign __DOLLAR__procmux__DOLLAR__654__A[12] = op_a[12];
  assign __DOLLAR__procmux__DOLLAR__654__A[13] = op_a[13];
  assign __DOLLAR__procmux__DOLLAR__654__A[14] = op_a[14];
  assign __DOLLAR__procmux__DOLLAR__654__A[15] = op_a[15];
  assign __DOLLAR__procmux__DOLLAR__654__A[2] = op_a[2];
  assign __DOLLAR__procmux__DOLLAR__654__A[3] = op_a[3];
  assign __DOLLAR__procmux__DOLLAR__654__A[4] = op_a[4];
  assign __DOLLAR__procmux__DOLLAR__654__A[5] = op_a[5];
  assign __DOLLAR__procmux__DOLLAR__654__A[6] = op_a[6];
  assign __DOLLAR__procmux__DOLLAR__654__A[7] = op_a[7];
  assign __DOLLAR__procmux__DOLLAR__654__A[8] = op_a[8];
  assign __DOLLAR__procmux__DOLLAR__654__A[9] = op_a[9];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__655_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__658_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__659_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__660_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__661_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__662_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__663_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__664_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__665_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__666_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__667_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__668_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__669_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__670_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__671_CMP0__A[5] = op_code[5];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[0] = op_code[0];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[1] = op_code[1];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[2] = op_code[2];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[3] = op_code[3];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[4] = op_code[4];
  assign __DOLLAR__procmux__DOLLAR__672_CMP0__A[5] = op_code[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[0] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[1] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[10] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[11] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[12] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[13] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[14] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[15] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[2] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[3] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[4] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[5] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[6] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[7] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[8] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__97__A[9] = __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__110__B[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__268__DOLLAR__109__Y[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[0] = op_b[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[1] = op_b[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[10] = op_b[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[11] = op_b[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[12] = op_b[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[13] = op_b[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[14] = op_b[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[15] = op_b[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[16] = op_a[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[17] = op_a[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[18] = op_a[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[19] = op_a[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[2] = op_b[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[20] = op_a[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[21] = op_a[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[22] = op_a[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[23] = op_a[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[24] = op_a[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[25] = op_a[9];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[26] = op_a[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[27] = op_a[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[28] = op_a[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[29] = op_a[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[3] = op_b[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[30] = op_a[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[31] = op_a[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[4] = op_b[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[5] = op_b[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[6] = op_b[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[7] = op_b[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[8] = op_b[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__122__A[9] = op_b[9];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[0] = test_mult_add__res[16];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[1] = test_mult_add__res[17];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[10] = test_mult_add__res[26];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[11] = test_mult_add__res[27];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[12] = test_mult_add__res[28];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[13] = test_mult_add__res[29];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[14] = test_mult_add__res[30];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[15] = test_mult_add__res[31];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[2] = test_mult_add__res[18];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[3] = test_mult_add__res[19];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[4] = test_mult_add__res[20];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[5] = test_mult_add__res[21];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[6] = test_mult_add__res[22];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[7] = test_mult_add__res[23];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[8] = test_mult_add__res[24];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__319__DOLLAR__125__A[9] = test_mult_add__res[25];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[0] = op_b[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[1] = op_b[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[10] = op_b[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[11] = op_b[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[12] = op_b[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[13] = op_b[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[14] = op_b[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[15] = op_b[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[16] = op_a[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[17] = op_a[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[18] = op_a[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[19] = op_a[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[2] = op_b[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[20] = op_a[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[21] = op_a[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[22] = op_a[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[23] = op_a[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[24] = op_a[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[25] = op_a[9];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[26] = op_a[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[27] = op_a[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[28] = op_a[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[29] = op_a[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[3] = op_b[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[30] = op_a[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[31] = op_a[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[4] = op_b[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[5] = op_b[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[6] = op_b[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[7] = op_b[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[8] = op_b[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__128__A[9] = op_b[9];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[0] = test_mult_add__res[24];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[1] = test_mult_add__res[25];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[2] = test_mult_add__res[26];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[3] = test_mult_add__res[27];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[4] = test_mult_add__res[28];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[5] = test_mult_add__res[29];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[6] = test_mult_add__res[30];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__330__DOLLAR__131__A[7] = test_mult_add__res[31];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[0] = op_a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[1] = op_a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[10] = op_a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[11] = op_a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[12] = op_a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[13] = op_a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[14] = op_a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[15] = op_a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[2] = op_a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[3] = op_a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[4] = op_a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[5] = op_a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[6] = op_a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[7] = op_a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[8] = op_a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__283__DOLLAR__114__B[9] = op_a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[0] = op_b[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[1] = op_b[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[10] = op_b[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[11] = op_b[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[12] = op_b[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[13] = op_b[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[14] = op_b[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[15] = op_b[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[2] = op_b[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[3] = op_b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[4] = op_b[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[5] = op_b[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[6] = op_b[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[7] = op_b[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[8] = op_b[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__A[9] = op_b[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[0] = op_a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[1] = op_a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[10] = op_a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[11] = op_a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[12] = op_a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[13] = op_a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[14] = op_a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[15] = op_a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[2] = op_a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[3] = op_a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[4] = op_a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[5] = op_a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[6] = op_a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[7] = op_a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[8] = op_a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__290__DOLLAR__116__B[9] = op_a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[0] = op_b[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[1] = op_b[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[10] = op_b[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[11] = op_b[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[12] = op_b[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[13] = op_b[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[14] = op_b[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[15] = op_b[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[2] = op_b[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[3] = op_b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[4] = op_b[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[5] = op_b[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[6] = op_b[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[7] = op_b[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[8] = op_b[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__A[9] = op_b[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[0] = op_a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[1] = op_a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[10] = op_a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[11] = op_a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[12] = op_a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[13] = op_a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[14] = op_a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[15] = op_a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[2] = op_a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[3] = op_a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[4] = op_a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[5] = op_a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[6] = op_a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[7] = op_a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[8] = op_a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__296__DOLLAR__118__B[9] = op_a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[0] = op_b[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[1] = op_b[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[10] = op_b[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[11] = op_b[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[12] = op_b[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[13] = op_b[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[14] = op_b[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[15] = op_b[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[2] = op_b[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[3] = op_b[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[4] = op_b[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[5] = op_b[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[6] = op_b[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[7] = op_b[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[8] = op_b[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__A[9] = op_b[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[0] = op_a[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[1] = op_a[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[10] = op_a[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[11] = op_a[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[12] = op_a[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[13] = op_a[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[14] = op_a[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[15] = op_a[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[2] = op_a[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[3] = op_a[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[4] = op_a[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[5] = op_a[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[6] = op_a[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[7] = op_a[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[8] = op_a[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__303__DOLLAR__119__B[9] = op_a[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__317__DOLLAR__124__B[0] = test_mult_add__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__328__DOLLAR__130__B[0] = test_mult_add__res[15];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[0] = op_a[0];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[1] = op_a[1];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[10] = op_a[10];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[11] = op_a[11];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[12] = op_a[12];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[13] = op_a[13];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[14] = op_a[14];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[15] = op_a[15];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[2] = op_a[2];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[3] = op_a[3];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[4] = op_a[4];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[5] = op_a[5];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[6] = op_a[6];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[7] = op_a[7];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[8] = op_a[8];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__A[9] = op_a[9];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[0] = op_b[0];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[1] = op_b[1];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[10] = op_b[10];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[11] = op_b[11];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[12] = op_b[12];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[13] = op_b[13];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[14] = op_b[14];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[15] = op_b[15];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[2] = op_b[2];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[3] = op_b[3];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[4] = op_b[4];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[5] = op_b[5];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[6] = op_b[6];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[7] = op_b[7];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[8] = op_b[8];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__181__DOLLAR__96__B[9] = op_b[9];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[0] = op_a[0];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[1] = op_a[1];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[10] = op_a[10];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[11] = op_a[11];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[12] = op_a[12];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[13] = op_a[13];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[14] = op_a[14];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[15] = op_a[15];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[2] = op_a[2];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[3] = op_a[3];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[4] = op_a[4];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[5] = op_a[5];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[6] = op_a[6];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[7] = op_a[7];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[8] = op_a[8];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__A[9] = op_a[9];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[0] = op_b[0];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[1] = op_b[1];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[10] = op_b[10];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[11] = op_b[11];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[12] = op_b[12];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[13] = op_b[13];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[14] = op_b[14];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[15] = op_b[15];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[2] = op_b[2];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[3] = op_b[3];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[4] = op_b[4];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[5] = op_b[5];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[6] = op_b[6];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[7] = op_b[7];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[8] = op_b[8];
  assign __DOLLAR__xor__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_comp_unq1__DOT__sv__COLON__347__DOLLAR__134__B[9] = op_b[9];
  assign test_mult_add__a[0] = op_a[0];
  assign test_shifter__a[0] = op_a[0];
  assign test_mult_add__a[1] = op_a[1];
  assign test_shifter__a[1] = op_a[1];
  assign test_mult_add__a[10] = op_a[10];
  assign test_shifter__a[10] = op_a[10];
  assign test_mult_add__a[11] = op_a[11];
  assign test_shifter__a[11] = op_a[11];
  assign test_mult_add__a[12] = op_a[12];
  assign test_shifter__a[12] = op_a[12];
  assign test_mult_add__a[13] = op_a[13];
  assign test_shifter__a[13] = op_a[13];
  assign test_mult_add__a[14] = op_a[14];
  assign test_shifter__a[14] = op_a[14];
  assign test_mult_add__a[15] = op_a[15];
  assign test_shifter__a[15] = op_a[15];
  assign test_mult_add__a[2] = op_a[2];
  assign test_shifter__a[2] = op_a[2];
  assign test_mult_add__a[3] = op_a[3];
  assign test_shifter__a[3] = op_a[3];
  assign test_mult_add__a[4] = op_a[4];
  assign test_shifter__a[4] = op_a[4];
  assign test_mult_add__a[5] = op_a[5];
  assign test_shifter__a[5] = op_a[5];
  assign test_mult_add__a[6] = op_a[6];
  assign test_shifter__a[6] = op_a[6];
  assign test_mult_add__a[7] = op_a[7];
  assign test_shifter__a[7] = op_a[7];
  assign test_mult_add__a[8] = op_a[8];
  assign test_shifter__a[8] = op_a[8];
  assign test_mult_add__a[9] = op_a[9];
  assign test_shifter__a[9] = op_a[9];
  assign test_mult_add__b[0] = op_b[0];
  assign test_shifter__b[0] = op_b[0];
  assign test_mult_add__b[1] = op_b[1];
  assign test_shifter__b[1] = op_b[1];
  assign test_mult_add__b[10] = op_b[10];
  assign test_mult_add__b[11] = op_b[11];
  assign test_mult_add__b[12] = op_b[12];
  assign test_mult_add__b[13] = op_b[13];
  assign test_mult_add__b[14] = op_b[14];
  assign test_mult_add__b[15] = op_b[15];
  assign test_mult_add__b[2] = op_b[2];
  assign test_shifter__b[2] = op_b[2];
  assign test_mult_add__b[3] = op_b[3];
  assign test_shifter__b[3] = op_b[3];
  assign test_mult_add__b[4] = op_b[4];
  assign test_mult_add__b[5] = op_b[5];
  assign test_mult_add__b[6] = op_b[6];
  assign test_mult_add__b[7] = op_b[7];
  assign test_mult_add__b[8] = op_b[8];
  assign test_mult_add__b[9] = op_b[9];

endmodule //test_pe_comp_unq1

module test_pe_unq1 (
  input  bit0,
  input  bit1,
  input  bit2,
  input [7:0] cfg_a,
  input [31:0] cfg_d,
  input  cfg_en,
  input  clk,
  input  clk_en,
  input [15:0] data0,
  input [15:0] data1,
  output  irq,
  output [15:0] read_data,
  output [15:0] res,
  output  res_p,
  input  rst_n
);
  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186' (Module and_U42)
  wire [1:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__A;
  wire [1:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__B;
  wire [1:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__Y;
  and_U42 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118' (Module reduce_or_U43)
  wire [9:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__Y;
  reduce_or_U43 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144' (Module reduce_or_U30)
  wire [3:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__Y;
  reduce_or_U30 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188' (Module reduce_or_U30)
  wire [3:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__Y;
  reduce_or_U30 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190' (Module rtMux_U8)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__S;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__Y;
  rtMux_U8 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176' (Module eq_U23)
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__A;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__Y;
  eq_U23 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163' (Module logic_not_U33)
  wire [0:0] __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__A;
  wire [0:0] __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y;
  logic_not_U33 __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163(
    .A(__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__A),
    .Y(__DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y)
  );

  //Wire declarations for instance '__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174' (Module ne_U34)
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__A;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__B;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__Y;
  ne_U34 __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174(
    .A(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__A),
    .B(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__B),
    .Y(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__Y)
  );

  //Wire declarations for instance '__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178' (Module ne_U34)
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__A;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__B;
  wire [0:0] __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__Y;
  ne_U34 __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178(
    .A(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__A),
    .B(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__B),
    .Y(__DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__Y)
  );

  //Wire declarations for instance '__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175' (Module not_U14)
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__A;
  wire [0:0] __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__Y;
  not_U14 __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175(
    .A(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__A),
    .Y(__DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__752' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__752__ARST;
  wire  __DOLLAR__procdff__DOLLAR__752__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__752__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__752__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__752(
    .ARST(__DOLLAR__procdff__DOLLAR__752__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__752__CLK),
    .D(__DOLLAR__procdff__DOLLAR__752__D),
    .Q(__DOLLAR__procdff__DOLLAR__752__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__753' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__753__ARST;
  wire  __DOLLAR__procdff__DOLLAR__753__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__753__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__753__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__753(
    .ARST(__DOLLAR__procdff__DOLLAR__753__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__753__CLK),
    .D(__DOLLAR__procdff__DOLLAR__753__D),
    .Q(__DOLLAR__procdff__DOLLAR__753__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__526_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__526_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__526_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__526_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__526_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__526_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__526_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__527_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__527_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__527_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__527_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__527_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__527_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__527_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__528_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__528_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__528_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__528_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__528_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__528_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__528_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__529_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__529_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__529_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__529_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__529_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__529_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__529_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__530_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__530_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__530_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__530_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__530_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__530_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__530_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__531_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__531_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__531_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__531_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__531_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__531_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__531_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__532_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__532_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__532_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__532_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__532_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__532_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__532_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__533_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__533_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__533_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__533_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__533_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__533_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__533_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__534_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__534_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__534_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__534_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__534_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__534_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__534_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__535_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__535_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__535_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__535_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__535_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__535_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__535_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__537_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__537_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__537_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__537_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__537_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__537_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__537_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__537_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__538_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__538_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__538_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__538_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__538_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__538_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__538_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__538_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__539_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__539_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__539_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__539_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__539_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__539_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__539_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__539_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__540_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__540_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__540_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__540_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__540_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__540_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__540_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__540_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__541_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__541_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__541_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__541_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__541_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__541_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__541_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__541_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__542_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__542_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__542_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__542_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__542_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__542_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__542_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__542_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__543_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__543_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__543_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__543_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__543_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__543_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__543_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__543_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__544_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__544_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__544_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__544_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__544_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__544_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__544_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__544_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__545_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__545_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__545_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__545_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__545_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__545_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__545_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__545_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__546_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__546_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__546_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__546_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__546_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__546_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__546_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__546_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__547_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__547_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__547_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__547_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__547_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__547_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__547_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__547_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__548_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__548_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__548_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__548_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__548_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__548_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__548_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__548_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__549_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__549_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__549_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__549_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__549_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__549_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__549_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__549_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__550_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__550_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__550_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__550_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__550_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__550_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__550_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__550_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__551_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__551_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__551_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__551_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__551_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__551_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__551_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__551_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__552_CMP0' (Module eq_U15)
  wire [3:0] __DOLLAR__procmux__DOLLAR__552_CMP0__A;
  wire [3:0] __DOLLAR__procmux__DOLLAR__552_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__552_CMP0__Y;
  eq_U15 __DOLLAR__procmux__DOLLAR__552_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__552_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__552_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__552_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__554' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__554__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__554__B;
  wire  __DOLLAR__procmux__DOLLAR__554__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__554__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__554(
    .A(__DOLLAR__procmux__DOLLAR__554__A),
    .B(__DOLLAR__procmux__DOLLAR__554__B),
    .S(__DOLLAR__procmux__DOLLAR__554__S),
    .Y(__DOLLAR__procmux__DOLLAR__554__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__557' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__557__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__557__B;
  wire  __DOLLAR__procmux__DOLLAR__557__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__557__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__557(
    .A(__DOLLAR__procmux__DOLLAR__557__A),
    .B(__DOLLAR__procmux__DOLLAR__557__B),
    .S(__DOLLAR__procmux__DOLLAR__557__S),
    .Y(__DOLLAR__procmux__DOLLAR__557__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143' (Module reduce_and_U44)
  wire [7:0] __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A;
  wire [0:0] __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__Y;
  reduce_and_U44 __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143(
    .A(__DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A),
    .Y(__DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162' (Module reduce_or_U37)
  wire [15:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__Y;
  reduce_or_U37 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__Y)
  );

  //Wire declarations for instance '__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187' (Module reduce_or_U13)
  wire [1:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__A;
  wire [0:0] __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__Y;
  reduce_or_U13 __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187(
    .A(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__A),
    .Y(__DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y)
  );

  //Wire declarations for instance 'test_debug_bit' (Module __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__1)
  wire  test_debug_bit__cfg_clk;
  wire  test_debug_bit__cfg_d;
  wire  test_debug_bit__cfg_en;
  wire  test_debug_bit__cfg_rst_n;
  wire  test_debug_bit__data_in;
  wire  test_debug_bit__debug_irq;
  __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__1 test_debug_bit(
    .cfg_clk(test_debug_bit__cfg_clk),
    .cfg_d(test_debug_bit__cfg_d),
    .cfg_en(test_debug_bit__cfg_en),
    .cfg_rst_n(test_debug_bit__cfg_rst_n),
    .data_in(test_debug_bit__data_in),
    .debug_irq(test_debug_bit__debug_irq)
  );

  //Wire declarations for instance 'test_debug_data' (Module __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__16)
  wire  test_debug_data__cfg_clk;
  wire [15:0] test_debug_data__cfg_d;
  wire  test_debug_data__cfg_en;
  wire  test_debug_data__cfg_rst_n;
  wire [15:0] test_debug_data__data_in;
  wire  test_debug_data__debug_irq;
  __DOLLAR__paramod__BACKSLASH__test_debug_reg__BACKSLASH__DataWidth__EQUALS__16 test_debug_data(
    .cfg_clk(test_debug_data__cfg_clk),
    .cfg_d(test_debug_data__cfg_d),
    .cfg_en(test_debug_data__cfg_en),
    .cfg_rst_n(test_debug_data__cfg_rst_n),
    .data_in(test_debug_data__data_in),
    .debug_irq(test_debug_data__debug_irq)
  );

  //Wire declarations for instance 'test_lut' (Module __DOLLAR__paramod__BACKSLASH__test_lut__BACKSLASH__DataWidth__EQUALS__1)
  wire [7:0] test_lut__cfg_a;
  wire  test_lut__cfg_clk;
  wire [31:0] test_lut__cfg_d;
  wire  test_lut__cfg_en;
  wire  test_lut__cfg_rst_n;
  wire  test_lut__op_a_in;
  wire  test_lut__op_b_in;
  wire  test_lut__op_c_in;
  wire  test_lut__res;
  __DOLLAR__paramod__BACKSLASH__test_lut__BACKSLASH__DataWidth__EQUALS__1 test_lut(
    .cfg_a(test_lut__cfg_a),
    .cfg_clk(test_lut__cfg_clk),
    .cfg_d(test_lut__cfg_d),
    .cfg_en(test_lut__cfg_en),
    .cfg_rst_n(test_lut__cfg_rst_n),
    .op_a_in(test_lut__op_a_in),
    .op_b_in(test_lut__op_b_in),
    .op_c_in(test_lut__op_c_in),
    .res(test_lut__res)
  );

  //Wire declarations for instance 'test_opt_reg_a' (Module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__16)
  wire  test_opt_reg_a__clk;
  wire  test_opt_reg_a__clk_en;
  wire [15:0] test_opt_reg_a__data_in;
  wire  test_opt_reg_a__load;
  wire [1:0] test_opt_reg_a__mode;
  wire [15:0] test_opt_reg_a__reg_data;
  wire [15:0] test_opt_reg_a__res;
  wire  test_opt_reg_a__rst_n;
  wire [15:0] test_opt_reg_a__val;
  __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__16 test_opt_reg_a(
    .clk(test_opt_reg_a__clk),
    .clk_en(test_opt_reg_a__clk_en),
    .data_in(test_opt_reg_a__data_in),
    .load(test_opt_reg_a__load),
    .mode(test_opt_reg_a__mode),
    .reg_data(test_opt_reg_a__reg_data),
    .res(test_opt_reg_a__res),
    .rst_n(test_opt_reg_a__rst_n),
    .val(test_opt_reg_a__val)
  );

  //Wire declarations for instance 'test_opt_reg_d' (Module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1)
  wire  test_opt_reg_d__clk;
  wire  test_opt_reg_d__clk_en;
  wire  test_opt_reg_d__data_in;
  wire  test_opt_reg_d__load;
  wire [1:0] test_opt_reg_d__mode;
  wire  test_opt_reg_d__reg_data;
  wire  test_opt_reg_d__res;
  wire  test_opt_reg_d__rst_n;
  wire  test_opt_reg_d__val;
  __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1 test_opt_reg_d(
    .clk(test_opt_reg_d__clk),
    .clk_en(test_opt_reg_d__clk_en),
    .data_in(test_opt_reg_d__data_in),
    .load(test_opt_reg_d__load),
    .mode(test_opt_reg_d__mode),
    .reg_data(test_opt_reg_d__reg_data),
    .res(test_opt_reg_d__res),
    .rst_n(test_opt_reg_d__rst_n),
    .val(test_opt_reg_d__val)
  );

  //Wire declarations for instance 'test_opt_reg_e' (Module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1)
  wire  test_opt_reg_e__clk;
  wire  test_opt_reg_e__clk_en;
  wire  test_opt_reg_e__data_in;
  wire  test_opt_reg_e__load;
  wire [1:0] test_opt_reg_e__mode;
  wire  test_opt_reg_e__reg_data;
  wire  test_opt_reg_e__res;
  wire  test_opt_reg_e__rst_n;
  wire  test_opt_reg_e__val;
  __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1 test_opt_reg_e(
    .clk(test_opt_reg_e__clk),
    .clk_en(test_opt_reg_e__clk_en),
    .data_in(test_opt_reg_e__data_in),
    .load(test_opt_reg_e__load),
    .mode(test_opt_reg_e__mode),
    .reg_data(test_opt_reg_e__reg_data),
    .res(test_opt_reg_e__res),
    .rst_n(test_opt_reg_e__rst_n),
    .val(test_opt_reg_e__val)
  );

  //Wire declarations for instance 'test_opt_reg_f' (Module __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1)
  wire  test_opt_reg_f__clk;
  wire  test_opt_reg_f__clk_en;
  wire  test_opt_reg_f__data_in;
  wire  test_opt_reg_f__load;
  wire [1:0] test_opt_reg_f__mode;
  wire  test_opt_reg_f__reg_data;
  wire  test_opt_reg_f__res;
  wire  test_opt_reg_f__rst_n;
  wire  test_opt_reg_f__val;
  __DOLLAR__paramod__BACKSLASH__test_opt_reg__BACKSLASH__DataWidth__EQUALS__1 test_opt_reg_f(
    .clk(test_opt_reg_f__clk),
    .clk_en(test_opt_reg_f__clk_en),
    .data_in(test_opt_reg_f__data_in),
    .load(test_opt_reg_f__load),
    .mode(test_opt_reg_f__mode),
    .reg_data(test_opt_reg_f__reg_data),
    .res(test_opt_reg_f__res),
    .rst_n(test_opt_reg_f__rst_n),
    .val(test_opt_reg_f__val)
  );

  //Wire declarations for instance 'test_opt_reg_file' (Module __DOLLAR__paramod__BACKSLASH__test_opt_reg_file__BACKSLASH__DataWidth__EQUALS__16)
  wire [7:0] test_opt_reg_file__cfg_a;
  wire [15:0] test_opt_reg_file__cfg_d;
  wire  test_opt_reg_file__cfg_en;
  wire  test_opt_reg_file__clk;
  wire  test_opt_reg_file__clk_en;
  wire [15:0] test_opt_reg_file__data_in;
  wire  test_opt_reg_file__load;
  wire [2:0] test_opt_reg_file__mode;
  wire [15:0] test_opt_reg_file__reg_data;
  wire [15:0] test_opt_reg_file__res;
  wire  test_opt_reg_file__rst_n;
  wire [15:0] test_opt_reg_file__val;
  __DOLLAR__paramod__BACKSLASH__test_opt_reg_file__BACKSLASH__DataWidth__EQUALS__16 test_opt_reg_file(
    .cfg_a(test_opt_reg_file__cfg_a),
    .cfg_d(test_opt_reg_file__cfg_d),
    .cfg_en(test_opt_reg_file__cfg_en),
    .clk(test_opt_reg_file__clk),
    .clk_en(test_opt_reg_file__clk_en),
    .data_in(test_opt_reg_file__data_in),
    .load(test_opt_reg_file__load),
    .mode(test_opt_reg_file__mode),
    .reg_data(test_opt_reg_file__reg_data),
    .res(test_opt_reg_file__res),
    .rst_n(test_opt_reg_file__rst_n),
    .val(test_opt_reg_file__val)
  );

  //Wire declarations for instance 'test_pe_comp' (Module test_pe_comp_unq1)
  wire  test_pe_comp__carry_out;
  wire [15:0] test_pe_comp__op_a;
  wire [15:0] test_pe_comp__op_b;
  wire [7:0] test_pe_comp__op_code;
  wire  test_pe_comp__op_d_p;
  wire  test_pe_comp__ovfl;
  wire [15:0] test_pe_comp__res;
  wire  test_pe_comp__res_p;
  test_pe_comp_unq1 test_pe_comp(
    .carry_out(test_pe_comp__carry_out),
    .op_a(test_pe_comp__op_a),
    .op_b(test_pe_comp__op_b),
    .op_code(test_pe_comp__op_code),
    .op_d_p(test_pe_comp__op_d_p),
    .ovfl(test_pe_comp__ovfl),
    .res(test_pe_comp__res),
    .res_p(test_pe_comp__res_p)
  );

  //All the connections
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__S = __DOLLAR__procmux__DOLLAR__526_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__S = __DOLLAR__procmux__DOLLAR__529_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__S = __DOLLAR__procmux__DOLLAR__528_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__S = __DOLLAR__procmux__DOLLAR__532_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__S = __DOLLAR__procmux__DOLLAR__531_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__S = __DOLLAR__procmux__DOLLAR__535_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__S = __DOLLAR__procmux__DOLLAR__534_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__S = __DOLLAR__procmux__DOLLAR__537_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__S = __DOLLAR__procmux__DOLLAR__539_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__S = __DOLLAR__procmux__DOLLAR__541_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__S = __DOLLAR__procmux__DOLLAR__543_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__S = __DOLLAR__procmux__DOLLAR__545_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__S = __DOLLAR__procmux__DOLLAR__547_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__S = __DOLLAR__procmux__DOLLAR__549_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__S = __DOLLAR__procmux__DOLLAR__551_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procdff__DOLLAR__752__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__752__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__753__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__753__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__526_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__527_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__528_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__529_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__530_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__531_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__532_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__533_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__534_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__535_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__537_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__538_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__539_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__540_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__541_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__542_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__543_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__544_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__545_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__546_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__547_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__548_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__549_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__550_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__551_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__552_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__554__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__Y[0];
  assign __DOLLAR__procmux__DOLLAR__557__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__S = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__S = __DOLLAR__procdff__DOLLAR__752__Q[9];
  assign test_opt_reg_d__data_in = bit0;
  assign test_opt_reg_e__data_in = bit1;
  assign test_opt_reg_f__data_in = bit2;
  assign test_lut__cfg_en = cfg_en;
  assign test_opt_reg_file__cfg_en = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__A[0] = cfg_en;
  assign test_debug_bit__cfg_clk = clk;
  assign test_debug_data__cfg_clk = clk;
  assign test_lut__cfg_clk = clk;
  assign test_opt_reg_a__clk = clk;
  assign test_opt_reg_d__clk = clk;
  assign test_opt_reg_e__clk = clk;
  assign test_opt_reg_f__clk = clk;
  assign test_opt_reg_file__clk = clk;
  assign test_opt_reg_a__clk_en = clk_en;
  assign test_opt_reg_d__clk_en = clk_en;
  assign test_opt_reg_e__clk_en = clk_en;
  assign test_opt_reg_f__clk_en = clk_en;
  assign test_opt_reg_file__clk_en = clk_en;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__A[0] = clk_en;
  assign irq = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__Y[0];
  assign res_p = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__Y[0];
  assign test_debug_bit__cfg_rst_n = rst_n;
  assign test_debug_data__cfg_rst_n = rst_n;
  assign test_lut__cfg_rst_n = rst_n;
  assign test_opt_reg_a__rst_n = rst_n;
  assign test_opt_reg_d__rst_n = rst_n;
  assign test_opt_reg_e__rst_n = rst_n;
  assign test_opt_reg_f__rst_n = rst_n;
  assign test_opt_reg_file__rst_n = rst_n;
  assign test_debug_bit__cfg_d = cfg_d[0];
  assign test_debug_bit__cfg_en = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__Y[0];
  assign test_debug_bit__data_in = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__A[0] = test_debug_bit__debug_irq;
  assign test_debug_data__cfg_en = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__A[1] = test_debug_data__debug_irq;
  assign test_lut__op_a_in = test_opt_reg_d__res;
  assign test_lut__op_b_in = test_opt_reg_e__res;
  assign test_lut__op_c_in = test_opt_reg_f__res;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__A[0] = test_lut__res;
  assign test_opt_reg_a__load = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__Y[0];
  assign test_opt_reg_d__load = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__A[0] = test_opt_reg_d__reg_data;
  assign test_pe_comp__op_d_p = test_opt_reg_d__res;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__B[0] = test_opt_reg_d__res;
  assign test_opt_reg_d__val = cfg_d[0];
  assign test_opt_reg_e__load = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__B[0] = test_opt_reg_e__reg_data;
  assign test_opt_reg_e__val = cfg_d[0];
  assign test_opt_reg_f__load = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__B[0] = test_opt_reg_f__reg_data;
  assign test_opt_reg_f__val = cfg_d[0];
  assign test_opt_reg_file__load = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__A[0] = test_pe_comp__carry_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__A[0] = test_pe_comp__carry_out;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__A[0] = test_pe_comp__carry_out;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__A[0] = test_pe_comp__carry_out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__A[0] = test_pe_comp__ovfl;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__B[0] = test_pe_comp__ovfl;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__B[0] = test_pe_comp__ovfl;
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__B[0] = test_pe_comp__ovfl;
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__B[0] = test_pe_comp__ovfl;
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__A[0] = test_pe_comp__ovfl;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__B[0] = test_pe_comp__res_p;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__B[0] = __DOLLAR__procdff__DOLLAR__752__Q[9];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__149__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__153__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[9];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__170__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__177__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__B[0] = __DOLLAR__procdff__DOLLAR__752__Q[10];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__B[1] = __DOLLAR__procdff__DOLLAR__752__Q[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__A[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__Y[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__187__A[1] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__417__DOLLAR__186__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[0] = __DOLLAR__procmux__DOLLAR__526_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[1] = __DOLLAR__procmux__DOLLAR__527_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[2] = __DOLLAR__procmux__DOLLAR__528_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[3] = __DOLLAR__procmux__DOLLAR__529_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[4] = __DOLLAR__procmux__DOLLAR__530_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[5] = __DOLLAR__procmux__DOLLAR__531_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[6] = __DOLLAR__procmux__DOLLAR__532_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[7] = __DOLLAR__procmux__DOLLAR__533_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[8] = __DOLLAR__procmux__DOLLAR__534_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__A[9] = __DOLLAR__procmux__DOLLAR__535_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__1120__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__1118__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__A[0] = __DOLLAR__procmux__DOLLAR__527_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__B[0] = __DOLLAR__procmux__DOLLAR__526_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1128__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__A[0] = __DOLLAR__procmux__DOLLAR__538_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__B[0] = __DOLLAR__procmux__DOLLAR__537_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1152__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__A[0] = __DOLLAR__procmux__DOLLAR__542_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__B[0] = __DOLLAR__procmux__DOLLAR__541_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1160__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__A[0] = __DOLLAR__procmux__DOLLAR__546_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__B[0] = __DOLLAR__procmux__DOLLAR__545_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1172__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__A[0] = __DOLLAR__procmux__DOLLAR__550_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__1180__B[0] = __DOLLAR__procmux__DOLLAR__549_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__A[0] = __DOLLAR__procmux__DOLLAR__533_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__A[1] = __DOLLAR__procmux__DOLLAR__532_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1140__A[2] = __DOLLAR__procmux__DOLLAR__531_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A[0] = __DOLLAR__procmux__DOLLAR__530_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A[1] = __DOLLAR__procmux__DOLLAR__529_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1144__A[2] = __DOLLAR__procmux__DOLLAR__528_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__A[0] = __DOLLAR__procmux__DOLLAR__540_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__A[1] = __DOLLAR__procmux__DOLLAR__539_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1164__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__A[0] = __DOLLAR__procmux__DOLLAR__548_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1184__A[1] = __DOLLAR__procmux__DOLLAR__547_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A[0] = __DOLLAR__procmux__DOLLAR__544_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__37__COLON__or_generator__DOLLAR__1188__A[1] = __DOLLAR__procmux__DOLLAR__543_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[0] = __DOLLAR__procdff__DOLLAR__753__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[1] = __DOLLAR__procdff__DOLLAR__753__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[10] = __DOLLAR__procdff__DOLLAR__753__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[11] = __DOLLAR__procdff__DOLLAR__753__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[12] = __DOLLAR__procdff__DOLLAR__753__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[13] = __DOLLAR__procdff__DOLLAR__753__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[14] = __DOLLAR__procdff__DOLLAR__753__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[15] = __DOLLAR__procdff__DOLLAR__753__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[2] = __DOLLAR__procdff__DOLLAR__753__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[3] = __DOLLAR__procdff__DOLLAR__753__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[4] = __DOLLAR__procdff__DOLLAR__753__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[5] = __DOLLAR__procdff__DOLLAR__753__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[6] = __DOLLAR__procdff__DOLLAR__753__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[7] = __DOLLAR__procdff__DOLLAR__753__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[8] = __DOLLAR__procdff__DOLLAR__753__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__A[9] = __DOLLAR__procdff__DOLLAR__753__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[0] = __DOLLAR__procdff__DOLLAR__752__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[1] = __DOLLAR__procdff__DOLLAR__752__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[10] = __DOLLAR__procdff__DOLLAR__752__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[11] = __DOLLAR__procdff__DOLLAR__752__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[12] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[13] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[14] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[15] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[2] = __DOLLAR__procdff__DOLLAR__752__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[3] = __DOLLAR__procdff__DOLLAR__752__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[4] = __DOLLAR__procdff__DOLLAR__752__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[5] = __DOLLAR__procdff__DOLLAR__752__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[6] = __DOLLAR__procdff__DOLLAR__752__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[7] = __DOLLAR__procdff__DOLLAR__752__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[8] = __DOLLAR__procdff__DOLLAR__752__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__B[9] = __DOLLAR__procdff__DOLLAR__752__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1122__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1124__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1126__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1130__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[0] = test_opt_reg_file__reg_data[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[1] = test_opt_reg_file__reg_data[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[10] = test_opt_reg_file__reg_data[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[11] = test_opt_reg_file__reg_data[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[12] = test_opt_reg_file__reg_data[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[13] = test_opt_reg_file__reg_data[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[14] = test_opt_reg_file__reg_data[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[15] = test_opt_reg_file__reg_data[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[2] = test_opt_reg_file__reg_data[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[3] = test_opt_reg_file__reg_data[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[4] = test_opt_reg_file__reg_data[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[5] = test_opt_reg_file__reg_data[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[6] = test_opt_reg_file__reg_data[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[7] = test_opt_reg_file__reg_data[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[8] = test_opt_reg_file__reg_data[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__A[9] = test_opt_reg_file__reg_data[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[0] = test_opt_reg_a__reg_data[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[1] = test_opt_reg_a__reg_data[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[10] = test_opt_reg_a__reg_data[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[11] = test_opt_reg_a__reg_data[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[12] = test_opt_reg_a__reg_data[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[13] = test_opt_reg_a__reg_data[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[14] = test_opt_reg_a__reg_data[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[15] = test_opt_reg_a__reg_data[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[2] = test_opt_reg_a__reg_data[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[3] = test_opt_reg_a__reg_data[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[4] = test_opt_reg_a__reg_data[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[5] = test_opt_reg_a__reg_data[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[6] = test_opt_reg_a__reg_data[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[7] = test_opt_reg_a__reg_data[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[8] = test_opt_reg_a__reg_data[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__B[9] = test_opt_reg_a__reg_data[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1132__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[0] = test_opt_reg_file__reg_data[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[1] = test_opt_reg_file__reg_data[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[10] = test_opt_reg_file__reg_data[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[11] = test_opt_reg_file__reg_data[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[12] = test_opt_reg_file__reg_data[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[13] = test_opt_reg_file__reg_data[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[14] = test_opt_reg_file__reg_data[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[15] = test_opt_reg_file__reg_data[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[2] = test_opt_reg_file__reg_data[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[3] = test_opt_reg_file__reg_data[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[4] = test_opt_reg_file__reg_data[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[5] = test_opt_reg_file__reg_data[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[6] = test_opt_reg_file__reg_data[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[7] = test_opt_reg_file__reg_data[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[8] = test_opt_reg_file__reg_data[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__B[9] = test_opt_reg_file__reg_data[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1134__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[0] = test_opt_reg_file__reg_data[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[1] = test_opt_reg_file__reg_data[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[10] = test_opt_reg_file__reg_data[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[11] = test_opt_reg_file__reg_data[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[12] = test_opt_reg_file__reg_data[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[13] = test_opt_reg_file__reg_data[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[14] = test_opt_reg_file__reg_data[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[15] = test_opt_reg_file__reg_data[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[2] = test_opt_reg_file__reg_data[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[3] = test_opt_reg_file__reg_data[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[4] = test_opt_reg_file__reg_data[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[5] = test_opt_reg_file__reg_data[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[6] = test_opt_reg_file__reg_data[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[7] = test_opt_reg_file__reg_data[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[8] = test_opt_reg_file__reg_data[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__B[9] = test_opt_reg_file__reg_data[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1136__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[0] = test_opt_reg_file__reg_data[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[1] = test_opt_reg_file__reg_data[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[10] = test_opt_reg_file__reg_data[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[11] = test_opt_reg_file__reg_data[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[12] = test_opt_reg_file__reg_data[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[13] = test_opt_reg_file__reg_data[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[14] = test_opt_reg_file__reg_data[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[15] = test_opt_reg_file__reg_data[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[2] = test_opt_reg_file__reg_data[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[3] = test_opt_reg_file__reg_data[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[4] = test_opt_reg_file__reg_data[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[5] = test_opt_reg_file__reg_data[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[6] = test_opt_reg_file__reg_data[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[7] = test_opt_reg_file__reg_data[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[8] = test_opt_reg_file__reg_data[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__B[9] = test_opt_reg_file__reg_data[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1138__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1142__Y[9];
  assign read_data[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[0];
  assign read_data[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[1];
  assign read_data[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[10];
  assign read_data[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[11];
  assign read_data[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[12];
  assign read_data[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[13];
  assign read_data[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[14];
  assign read_data[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[15];
  assign read_data[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[2];
  assign read_data[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[3];
  assign read_data[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[4];
  assign read_data[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[5];
  assign read_data[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[6];
  assign read_data[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[7];
  assign read_data[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[8];
  assign read_data[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1146__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1148__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__B[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1150__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1154__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__B[0] = __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1156__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__B[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1158__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1162__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1166__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__339__DOLLAR__168__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1168__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1170__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1174__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__335__DOLLAR__166__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1176__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__B[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1178__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1182__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1190__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__1186__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__146__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__177__DOLLAR__145__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__147__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__152__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__198__DOLLAR__151__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__157__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__230__DOLLAR__156__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__159__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__244__DOLLAR__158__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__161__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__259__DOLLAR__160__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__342__DOLLAR__173__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__176__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__183__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__395__DOLLAR__182__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__185__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__407__DOLLAR__184__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__144__B[0] = __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__150__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__197__DOLLAR__148__Y[0];
  assign __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__A[0] = __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__333__DOLLAR__165__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__340__DOLLAR__169__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__344__DOLLAR__175__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__B[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__A[0] = __DOLLAR__logic_not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__163__Y[0];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__343__DOLLAR__174__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__179__B[0] = __DOLLAR__ne__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__345__DOLLAR__178__Y[0];
  assign __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__337__DOLLAR__167__A[0] = test_pe_comp__res[15];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__172__A[0] = __DOLLAR__not__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__341__DOLLAR__171__Y[0];
  assign __DOLLAR__procdff__DOLLAR__752__D[0] = __DOLLAR__procmux__DOLLAR__557__Y[0];
  assign __DOLLAR__procdff__DOLLAR__752__D[1] = __DOLLAR__procmux__DOLLAR__557__Y[1];
  assign __DOLLAR__procdff__DOLLAR__752__D[10] = __DOLLAR__procmux__DOLLAR__557__Y[10];
  assign __DOLLAR__procdff__DOLLAR__752__D[11] = __DOLLAR__procmux__DOLLAR__557__Y[11];
  assign __DOLLAR__procdff__DOLLAR__752__D[12] = __DOLLAR__procmux__DOLLAR__557__Y[12];
  assign __DOLLAR__procdff__DOLLAR__752__D[13] = __DOLLAR__procmux__DOLLAR__557__Y[13];
  assign __DOLLAR__procdff__DOLLAR__752__D[14] = __DOLLAR__procmux__DOLLAR__557__Y[14];
  assign __DOLLAR__procdff__DOLLAR__752__D[15] = __DOLLAR__procmux__DOLLAR__557__Y[15];
  assign __DOLLAR__procdff__DOLLAR__752__D[2] = __DOLLAR__procmux__DOLLAR__557__Y[2];
  assign __DOLLAR__procdff__DOLLAR__752__D[3] = __DOLLAR__procmux__DOLLAR__557__Y[3];
  assign __DOLLAR__procdff__DOLLAR__752__D[4] = __DOLLAR__procmux__DOLLAR__557__Y[4];
  assign __DOLLAR__procdff__DOLLAR__752__D[5] = __DOLLAR__procmux__DOLLAR__557__Y[5];
  assign __DOLLAR__procdff__DOLLAR__752__D[6] = __DOLLAR__procmux__DOLLAR__557__Y[6];
  assign __DOLLAR__procdff__DOLLAR__752__D[7] = __DOLLAR__procmux__DOLLAR__557__Y[7];
  assign __DOLLAR__procdff__DOLLAR__752__D[8] = __DOLLAR__procmux__DOLLAR__557__Y[8];
  assign __DOLLAR__procdff__DOLLAR__752__D[9] = __DOLLAR__procmux__DOLLAR__557__Y[9];
  assign __DOLLAR__procmux__DOLLAR__557__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[0];
  assign test_pe_comp__op_code[0] = __DOLLAR__procdff__DOLLAR__752__Q[0];
  assign __DOLLAR__procmux__DOLLAR__557__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[1];
  assign test_pe_comp__op_code[1] = __DOLLAR__procdff__DOLLAR__752__Q[1];
  assign __DOLLAR__procmux__DOLLAR__557__A[10] = __DOLLAR__procdff__DOLLAR__752__Q[10];
  assign __DOLLAR__procmux__DOLLAR__557__A[11] = __DOLLAR__procdff__DOLLAR__752__Q[11];
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__A[0] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__557__A[12] = __DOLLAR__procdff__DOLLAR__752__Q[12];
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__A[1] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__557__A[13] = __DOLLAR__procdff__DOLLAR__752__Q[13];
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__557__A[14] = __DOLLAR__procdff__DOLLAR__752__Q[14];
  assign __DOLLAR__procmux__DOLLAR__537_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__538_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__539_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__540_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__541_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__542_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__543_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__544_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__545_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__546_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__547_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__548_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__549_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__550_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__551_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__552_CMP0__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__557__A[15] = __DOLLAR__procdff__DOLLAR__752__Q[15];
  assign __DOLLAR__procmux__DOLLAR__557__A[2] = __DOLLAR__procdff__DOLLAR__752__Q[2];
  assign test_pe_comp__op_code[2] = __DOLLAR__procdff__DOLLAR__752__Q[2];
  assign __DOLLAR__procmux__DOLLAR__557__A[3] = __DOLLAR__procdff__DOLLAR__752__Q[3];
  assign test_pe_comp__op_code[3] = __DOLLAR__procdff__DOLLAR__752__Q[3];
  assign __DOLLAR__procmux__DOLLAR__557__A[4] = __DOLLAR__procdff__DOLLAR__752__Q[4];
  assign test_pe_comp__op_code[4] = __DOLLAR__procdff__DOLLAR__752__Q[4];
  assign __DOLLAR__procmux__DOLLAR__557__A[5] = __DOLLAR__procdff__DOLLAR__752__Q[5];
  assign test_pe_comp__op_code[5] = __DOLLAR__procdff__DOLLAR__752__Q[5];
  assign __DOLLAR__procmux__DOLLAR__557__A[6] = __DOLLAR__procdff__DOLLAR__752__Q[6];
  assign test_pe_comp__op_code[6] = __DOLLAR__procdff__DOLLAR__752__Q[6];
  assign __DOLLAR__procmux__DOLLAR__557__A[7] = __DOLLAR__procdff__DOLLAR__752__Q[7];
  assign test_pe_comp__op_code[7] = __DOLLAR__procdff__DOLLAR__752__Q[7];
  assign __DOLLAR__procmux__DOLLAR__557__A[8] = __DOLLAR__procdff__DOLLAR__752__Q[8];
  assign __DOLLAR__procmux__DOLLAR__557__A[9] = __DOLLAR__procdff__DOLLAR__752__Q[9];
  assign __DOLLAR__procdff__DOLLAR__753__D[0] = __DOLLAR__procmux__DOLLAR__554__Y[0];
  assign __DOLLAR__procdff__DOLLAR__753__D[1] = __DOLLAR__procmux__DOLLAR__554__Y[1];
  assign __DOLLAR__procdff__DOLLAR__753__D[10] = __DOLLAR__procmux__DOLLAR__554__Y[10];
  assign __DOLLAR__procdff__DOLLAR__753__D[11] = __DOLLAR__procmux__DOLLAR__554__Y[11];
  assign __DOLLAR__procdff__DOLLAR__753__D[12] = __DOLLAR__procmux__DOLLAR__554__Y[12];
  assign __DOLLAR__procdff__DOLLAR__753__D[13] = __DOLLAR__procmux__DOLLAR__554__Y[13];
  assign __DOLLAR__procdff__DOLLAR__753__D[14] = __DOLLAR__procmux__DOLLAR__554__Y[14];
  assign __DOLLAR__procdff__DOLLAR__753__D[15] = __DOLLAR__procmux__DOLLAR__554__Y[15];
  assign __DOLLAR__procdff__DOLLAR__753__D[2] = __DOLLAR__procmux__DOLLAR__554__Y[2];
  assign __DOLLAR__procdff__DOLLAR__753__D[3] = __DOLLAR__procmux__DOLLAR__554__Y[3];
  assign __DOLLAR__procdff__DOLLAR__753__D[4] = __DOLLAR__procmux__DOLLAR__554__Y[4];
  assign __DOLLAR__procdff__DOLLAR__753__D[5] = __DOLLAR__procmux__DOLLAR__554__Y[5];
  assign __DOLLAR__procdff__DOLLAR__753__D[6] = __DOLLAR__procmux__DOLLAR__554__Y[6];
  assign __DOLLAR__procdff__DOLLAR__753__D[7] = __DOLLAR__procmux__DOLLAR__554__Y[7];
  assign __DOLLAR__procdff__DOLLAR__753__D[8] = __DOLLAR__procmux__DOLLAR__554__Y[8];
  assign __DOLLAR__procdff__DOLLAR__753__D[9] = __DOLLAR__procmux__DOLLAR__554__Y[9];
  assign __DOLLAR__procmux__DOLLAR__554__A[0] = __DOLLAR__procdff__DOLLAR__753__Q[0];
  assign test_opt_reg_a__mode[0] = __DOLLAR__procdff__DOLLAR__753__Q[0];
  assign __DOLLAR__procmux__DOLLAR__554__A[1] = __DOLLAR__procdff__DOLLAR__753__Q[1];
  assign test_opt_reg_a__mode[1] = __DOLLAR__procdff__DOLLAR__753__Q[1];
  assign __DOLLAR__procmux__DOLLAR__554__A[10] = __DOLLAR__procdff__DOLLAR__753__Q[10];
  assign test_opt_reg_e__mode[0] = __DOLLAR__procdff__DOLLAR__753__Q[10];
  assign __DOLLAR__procmux__DOLLAR__554__A[11] = __DOLLAR__procdff__DOLLAR__753__Q[11];
  assign test_opt_reg_e__mode[1] = __DOLLAR__procdff__DOLLAR__753__Q[11];
  assign __DOLLAR__procmux__DOLLAR__554__A[12] = __DOLLAR__procdff__DOLLAR__753__Q[12];
  assign test_opt_reg_f__mode[0] = __DOLLAR__procdff__DOLLAR__753__Q[12];
  assign __DOLLAR__procmux__DOLLAR__554__A[13] = __DOLLAR__procdff__DOLLAR__753__Q[13];
  assign test_opt_reg_f__mode[1] = __DOLLAR__procdff__DOLLAR__753__Q[13];
  assign __DOLLAR__procmux__DOLLAR__554__A[14] = __DOLLAR__procdff__DOLLAR__753__Q[14];
  assign __DOLLAR__procmux__DOLLAR__554__A[15] = __DOLLAR__procdff__DOLLAR__753__Q[15];
  assign __DOLLAR__procmux__DOLLAR__554__A[2] = __DOLLAR__procdff__DOLLAR__753__Q[2];
  assign test_opt_reg_file__mode[0] = __DOLLAR__procdff__DOLLAR__753__Q[2];
  assign __DOLLAR__procmux__DOLLAR__554__A[3] = __DOLLAR__procdff__DOLLAR__753__Q[3];
  assign test_opt_reg_file__mode[1] = __DOLLAR__procdff__DOLLAR__753__Q[3];
  assign __DOLLAR__procmux__DOLLAR__554__A[4] = __DOLLAR__procdff__DOLLAR__753__Q[4];
  assign test_opt_reg_file__mode[2] = __DOLLAR__procdff__DOLLAR__753__Q[4];
  assign __DOLLAR__procmux__DOLLAR__554__A[5] = __DOLLAR__procdff__DOLLAR__753__Q[5];
  assign __DOLLAR__procmux__DOLLAR__554__A[6] = __DOLLAR__procdff__DOLLAR__753__Q[6];
  assign __DOLLAR__procmux__DOLLAR__554__A[7] = __DOLLAR__procdff__DOLLAR__753__Q[7];
  assign __DOLLAR__procmux__DOLLAR__554__A[8] = __DOLLAR__procdff__DOLLAR__753__Q[8];
  assign test_opt_reg_d__mode[0] = __DOLLAR__procdff__DOLLAR__753__Q[8];
  assign __DOLLAR__procmux__DOLLAR__554__A[9] = __DOLLAR__procdff__DOLLAR__753__Q[9];
  assign test_opt_reg_d__mode[1] = __DOLLAR__procdff__DOLLAR__753__Q[9];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__526_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__527_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__528_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__529_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__530_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__531_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__532_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__533_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__534_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__535_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__554__B[0] = cfg_d[16];
  assign __DOLLAR__procmux__DOLLAR__554__B[1] = cfg_d[17];
  assign __DOLLAR__procmux__DOLLAR__554__B[10] = cfg_d[26];
  assign __DOLLAR__procmux__DOLLAR__554__B[11] = cfg_d[27];
  assign __DOLLAR__procmux__DOLLAR__554__B[12] = cfg_d[28];
  assign __DOLLAR__procmux__DOLLAR__554__B[13] = cfg_d[29];
  assign __DOLLAR__procmux__DOLLAR__554__B[14] = cfg_d[30];
  assign __DOLLAR__procmux__DOLLAR__554__B[15] = cfg_d[31];
  assign __DOLLAR__procmux__DOLLAR__554__B[2] = cfg_d[18];
  assign __DOLLAR__procmux__DOLLAR__554__B[3] = cfg_d[19];
  assign __DOLLAR__procmux__DOLLAR__554__B[4] = cfg_d[20];
  assign __DOLLAR__procmux__DOLLAR__554__B[5] = cfg_d[21];
  assign __DOLLAR__procmux__DOLLAR__554__B[6] = cfg_d[22];
  assign __DOLLAR__procmux__DOLLAR__554__B[7] = cfg_d[23];
  assign __DOLLAR__procmux__DOLLAR__554__B[8] = cfg_d[24];
  assign __DOLLAR__procmux__DOLLAR__554__B[9] = cfg_d[25];
  assign __DOLLAR__procmux__DOLLAR__557__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__557__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__557__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__557__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__557__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__557__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__557__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__557__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__557__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__557__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__557__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__557__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__557__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__557__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__557__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__557__B[9] = cfg_d[9];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[0] = cfg_a[0];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[1] = cfg_a[1];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[2] = cfg_a[2];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[3] = cfg_a[3];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[4] = cfg_a[4];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[5] = cfg_a[5];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[6] = cfg_a[6];
  assign __DOLLAR__reduce_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__160__DOLLAR__143__A[7] = cfg_a[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[0] = test_pe_comp__res[0];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[1] = test_pe_comp__res[1];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[10] = test_pe_comp__res[10];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[11] = test_pe_comp__res[11];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[12] = test_pe_comp__res[12];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[13] = test_pe_comp__res[13];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[14] = test_pe_comp__res[14];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[15] = test_pe_comp__res[15];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[2] = test_pe_comp__res[2];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[3] = test_pe_comp__res[3];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[4] = test_pe_comp__res[4];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[5] = test_pe_comp__res[5];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[6] = test_pe_comp__res[6];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[7] = test_pe_comp__res[7];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[8] = test_pe_comp__res[8];
  assign __DOLLAR__reduce_or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__309__DOLLAR__162__A[9] = test_pe_comp__res[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[0] = test_pe_comp__res[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[1] = test_pe_comp__res[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[10] = test_pe_comp__res[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[11] = test_pe_comp__res[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[12] = test_pe_comp__res[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[13] = test_pe_comp__res[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[14] = test_pe_comp__res[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[15] = test_pe_comp__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[2] = test_pe_comp__res[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[3] = test_pe_comp__res[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[4] = test_pe_comp__res[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[5] = test_pe_comp__res[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[6] = test_pe_comp__res[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[7] = test_pe_comp__res[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[8] = test_pe_comp__res[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__A[9] = test_pe_comp__res[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__A[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__154__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[0] = cfg_d[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[1] = cfg_d[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[10] = cfg_d[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[11] = cfg_d[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[12] = cfg_d[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[13] = cfg_d[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[14] = cfg_d[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[15] = cfg_d[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[2] = cfg_d[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[3] = cfg_d[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[4] = cfg_d[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[5] = cfg_d[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[6] = cfg_d[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[7] = cfg_d[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[8] = cfg_d[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__B[9] = cfg_d[9];
  assign test_opt_reg_file__val[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[0];
  assign test_opt_reg_file__val[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[1];
  assign test_opt_reg_file__val[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[10];
  assign test_opt_reg_file__val[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[11];
  assign test_opt_reg_file__val[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[12];
  assign test_opt_reg_file__val[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[13];
  assign test_opt_reg_file__val[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[14];
  assign test_opt_reg_file__val[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[15];
  assign test_opt_reg_file__val[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[2];
  assign test_opt_reg_file__val[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[3];
  assign test_opt_reg_file__val[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[4];
  assign test_opt_reg_file__val[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[5];
  assign test_opt_reg_file__val[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[6];
  assign test_opt_reg_file__val[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[7];
  assign test_opt_reg_file__val[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[8];
  assign test_opt_reg_file__val[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__200__DOLLAR__155__Y[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[0] = test_pe_comp__res[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[1] = test_pe_comp__res[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[10] = test_pe_comp__res[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[11] = test_pe_comp__res[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[12] = test_pe_comp__res[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[13] = test_pe_comp__res[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[14] = test_pe_comp__res[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[15] = test_pe_comp__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[2] = test_pe_comp__res[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[3] = test_pe_comp__res[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[4] = test_pe_comp__res[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[5] = test_pe_comp__res[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[6] = test_pe_comp__res[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[7] = test_pe_comp__res[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[8] = test_pe_comp__res[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__A[9] = test_pe_comp__res[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[0] = test_opt_reg_file__res[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[1] = test_opt_reg_file__res[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[10] = test_opt_reg_file__res[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[11] = test_opt_reg_file__res[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[12] = test_opt_reg_file__res[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[13] = test_opt_reg_file__res[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[14] = test_opt_reg_file__res[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[15] = test_opt_reg_file__res[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[2] = test_opt_reg_file__res[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[3] = test_opt_reg_file__res[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[4] = test_opt_reg_file__res[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[5] = test_opt_reg_file__res[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[6] = test_opt_reg_file__res[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[7] = test_opt_reg_file__res[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[8] = test_opt_reg_file__res[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__B[9] = test_opt_reg_file__res[9];
  assign res[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[0];
  assign test_debug_data__data_in[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[0];
  assign res[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[1];
  assign test_debug_data__data_in[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[1];
  assign res[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[10];
  assign test_debug_data__data_in[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[10];
  assign res[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[11];
  assign test_debug_data__data_in[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[11];
  assign res[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[12];
  assign test_debug_data__data_in[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[12];
  assign res[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[13];
  assign test_debug_data__data_in[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[13];
  assign res[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[14];
  assign test_debug_data__data_in[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[14];
  assign res[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[15];
  assign test_debug_data__data_in[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[15];
  assign res[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[2];
  assign test_debug_data__data_in[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[2];
  assign res[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[3];
  assign test_debug_data__data_in[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[3];
  assign res[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[4];
  assign test_debug_data__data_in[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[4];
  assign res[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[5];
  assign test_debug_data__data_in[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[5];
  assign res[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[6];
  assign test_debug_data__data_in[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[6];
  assign res[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[7];
  assign test_debug_data__data_in[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[7];
  assign res[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[8];
  assign test_debug_data__data_in[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[8];
  assign res[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[9];
  assign test_debug_data__data_in[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_pe_unq1__DOT__sv__COLON__380__DOLLAR__180__Y[9];
  assign test_lut__cfg_a[0] = cfg_a[0];
  assign test_opt_reg_file__cfg_a[0] = cfg_a[0];
  assign test_lut__cfg_a[1] = cfg_a[1];
  assign test_opt_reg_file__cfg_a[1] = cfg_a[1];
  assign test_lut__cfg_a[2] = cfg_a[2];
  assign test_opt_reg_file__cfg_a[2] = cfg_a[2];
  assign test_lut__cfg_a[3] = cfg_a[3];
  assign test_opt_reg_file__cfg_a[3] = cfg_a[3];
  assign test_lut__cfg_a[4] = cfg_a[4];
  assign test_opt_reg_file__cfg_a[4] = cfg_a[4];
  assign test_lut__cfg_a[5] = cfg_a[5];
  assign test_opt_reg_file__cfg_a[5] = cfg_a[5];
  assign test_lut__cfg_a[6] = cfg_a[6];
  assign test_opt_reg_file__cfg_a[6] = cfg_a[6];
  assign test_lut__cfg_a[7] = cfg_a[7];
  assign test_opt_reg_file__cfg_a[7] = cfg_a[7];
  assign test_debug_data__cfg_d[0] = cfg_d[0];
  assign test_lut__cfg_d[0] = cfg_d[0];
  assign test_opt_reg_a__val[0] = cfg_d[0];
  assign test_opt_reg_file__cfg_d[0] = cfg_d[0];
  assign test_debug_data__cfg_d[1] = cfg_d[1];
  assign test_lut__cfg_d[1] = cfg_d[1];
  assign test_opt_reg_a__val[1] = cfg_d[1];
  assign test_opt_reg_file__cfg_d[1] = cfg_d[1];
  assign test_debug_data__cfg_d[10] = cfg_d[10];
  assign test_lut__cfg_d[10] = cfg_d[10];
  assign test_opt_reg_a__val[10] = cfg_d[10];
  assign test_opt_reg_file__cfg_d[10] = cfg_d[10];
  assign test_debug_data__cfg_d[11] = cfg_d[11];
  assign test_lut__cfg_d[11] = cfg_d[11];
  assign test_opt_reg_a__val[11] = cfg_d[11];
  assign test_opt_reg_file__cfg_d[11] = cfg_d[11];
  assign test_debug_data__cfg_d[12] = cfg_d[12];
  assign test_lut__cfg_d[12] = cfg_d[12];
  assign test_opt_reg_a__val[12] = cfg_d[12];
  assign test_opt_reg_file__cfg_d[12] = cfg_d[12];
  assign test_debug_data__cfg_d[13] = cfg_d[13];
  assign test_lut__cfg_d[13] = cfg_d[13];
  assign test_opt_reg_a__val[13] = cfg_d[13];
  assign test_opt_reg_file__cfg_d[13] = cfg_d[13];
  assign test_debug_data__cfg_d[14] = cfg_d[14];
  assign test_lut__cfg_d[14] = cfg_d[14];
  assign test_opt_reg_a__val[14] = cfg_d[14];
  assign test_opt_reg_file__cfg_d[14] = cfg_d[14];
  assign test_debug_data__cfg_d[15] = cfg_d[15];
  assign test_lut__cfg_d[15] = cfg_d[15];
  assign test_opt_reg_a__val[15] = cfg_d[15];
  assign test_opt_reg_file__cfg_d[15] = cfg_d[15];
  assign test_lut__cfg_d[16] = cfg_d[16];
  assign test_lut__cfg_d[17] = cfg_d[17];
  assign test_lut__cfg_d[18] = cfg_d[18];
  assign test_lut__cfg_d[19] = cfg_d[19];
  assign test_debug_data__cfg_d[2] = cfg_d[2];
  assign test_lut__cfg_d[2] = cfg_d[2];
  assign test_opt_reg_a__val[2] = cfg_d[2];
  assign test_opt_reg_file__cfg_d[2] = cfg_d[2];
  assign test_lut__cfg_d[20] = cfg_d[20];
  assign test_lut__cfg_d[21] = cfg_d[21];
  assign test_lut__cfg_d[22] = cfg_d[22];
  assign test_lut__cfg_d[23] = cfg_d[23];
  assign test_lut__cfg_d[24] = cfg_d[24];
  assign test_lut__cfg_d[25] = cfg_d[25];
  assign test_lut__cfg_d[26] = cfg_d[26];
  assign test_lut__cfg_d[27] = cfg_d[27];
  assign test_lut__cfg_d[28] = cfg_d[28];
  assign test_lut__cfg_d[29] = cfg_d[29];
  assign test_debug_data__cfg_d[3] = cfg_d[3];
  assign test_lut__cfg_d[3] = cfg_d[3];
  assign test_opt_reg_a__val[3] = cfg_d[3];
  assign test_opt_reg_file__cfg_d[3] = cfg_d[3];
  assign test_lut__cfg_d[30] = cfg_d[30];
  assign test_lut__cfg_d[31] = cfg_d[31];
  assign test_debug_data__cfg_d[4] = cfg_d[4];
  assign test_lut__cfg_d[4] = cfg_d[4];
  assign test_opt_reg_a__val[4] = cfg_d[4];
  assign test_opt_reg_file__cfg_d[4] = cfg_d[4];
  assign test_debug_data__cfg_d[5] = cfg_d[5];
  assign test_lut__cfg_d[5] = cfg_d[5];
  assign test_opt_reg_a__val[5] = cfg_d[5];
  assign test_opt_reg_file__cfg_d[5] = cfg_d[5];
  assign test_debug_data__cfg_d[6] = cfg_d[6];
  assign test_lut__cfg_d[6] = cfg_d[6];
  assign test_opt_reg_a__val[6] = cfg_d[6];
  assign test_opt_reg_file__cfg_d[6] = cfg_d[6];
  assign test_debug_data__cfg_d[7] = cfg_d[7];
  assign test_lut__cfg_d[7] = cfg_d[7];
  assign test_opt_reg_a__val[7] = cfg_d[7];
  assign test_opt_reg_file__cfg_d[7] = cfg_d[7];
  assign test_debug_data__cfg_d[8] = cfg_d[8];
  assign test_lut__cfg_d[8] = cfg_d[8];
  assign test_opt_reg_a__val[8] = cfg_d[8];
  assign test_opt_reg_file__cfg_d[8] = cfg_d[8];
  assign test_debug_data__cfg_d[9] = cfg_d[9];
  assign test_lut__cfg_d[9] = cfg_d[9];
  assign test_opt_reg_a__val[9] = cfg_d[9];
  assign test_opt_reg_file__cfg_d[9] = cfg_d[9];
  assign test_opt_reg_a__data_in[0] = data0[0];
  assign test_opt_reg_a__data_in[1] = data0[1];
  assign test_opt_reg_a__data_in[10] = data0[10];
  assign test_opt_reg_a__data_in[11] = data0[11];
  assign test_opt_reg_a__data_in[12] = data0[12];
  assign test_opt_reg_a__data_in[13] = data0[13];
  assign test_opt_reg_a__data_in[14] = data0[14];
  assign test_opt_reg_a__data_in[15] = data0[15];
  assign test_opt_reg_a__data_in[2] = data0[2];
  assign test_opt_reg_a__data_in[3] = data0[3];
  assign test_opt_reg_a__data_in[4] = data0[4];
  assign test_opt_reg_a__data_in[5] = data0[5];
  assign test_opt_reg_a__data_in[6] = data0[6];
  assign test_opt_reg_a__data_in[7] = data0[7];
  assign test_opt_reg_a__data_in[8] = data0[8];
  assign test_opt_reg_a__data_in[9] = data0[9];
  assign test_opt_reg_file__data_in[0] = data1[0];
  assign test_opt_reg_file__data_in[1] = data1[1];
  assign test_opt_reg_file__data_in[10] = data1[10];
  assign test_opt_reg_file__data_in[11] = data1[11];
  assign test_opt_reg_file__data_in[12] = data1[12];
  assign test_opt_reg_file__data_in[13] = data1[13];
  assign test_opt_reg_file__data_in[14] = data1[14];
  assign test_opt_reg_file__data_in[15] = data1[15];
  assign test_opt_reg_file__data_in[2] = data1[2];
  assign test_opt_reg_file__data_in[3] = data1[3];
  assign test_opt_reg_file__data_in[4] = data1[4];
  assign test_opt_reg_file__data_in[5] = data1[5];
  assign test_opt_reg_file__data_in[6] = data1[6];
  assign test_opt_reg_file__data_in[7] = data1[7];
  assign test_opt_reg_file__data_in[8] = data1[8];
  assign test_opt_reg_file__data_in[9] = data1[9];
  assign test_pe_comp__op_a[0] = test_opt_reg_a__res[0];
  assign test_pe_comp__op_a[1] = test_opt_reg_a__res[1];
  assign test_pe_comp__op_a[10] = test_opt_reg_a__res[10];
  assign test_pe_comp__op_a[11] = test_opt_reg_a__res[11];
  assign test_pe_comp__op_a[12] = test_opt_reg_a__res[12];
  assign test_pe_comp__op_a[13] = test_opt_reg_a__res[13];
  assign test_pe_comp__op_a[14] = test_opt_reg_a__res[14];
  assign test_pe_comp__op_a[15] = test_opt_reg_a__res[15];
  assign test_pe_comp__op_a[2] = test_opt_reg_a__res[2];
  assign test_pe_comp__op_a[3] = test_opt_reg_a__res[3];
  assign test_pe_comp__op_a[4] = test_opt_reg_a__res[4];
  assign test_pe_comp__op_a[5] = test_opt_reg_a__res[5];
  assign test_pe_comp__op_a[6] = test_opt_reg_a__res[6];
  assign test_pe_comp__op_a[7] = test_opt_reg_a__res[7];
  assign test_pe_comp__op_a[8] = test_opt_reg_a__res[8];
  assign test_pe_comp__op_a[9] = test_opt_reg_a__res[9];
  assign test_pe_comp__op_b[0] = test_opt_reg_file__res[0];
  assign test_pe_comp__op_b[1] = test_opt_reg_file__res[1];
  assign test_pe_comp__op_b[10] = test_opt_reg_file__res[10];
  assign test_pe_comp__op_b[11] = test_opt_reg_file__res[11];
  assign test_pe_comp__op_b[12] = test_opt_reg_file__res[12];
  assign test_pe_comp__op_b[13] = test_opt_reg_file__res[13];
  assign test_pe_comp__op_b[14] = test_opt_reg_file__res[14];
  assign test_pe_comp__op_b[15] = test_opt_reg_file__res[15];
  assign test_pe_comp__op_b[2] = test_opt_reg_file__res[2];
  assign test_pe_comp__op_b[3] = test_opt_reg_file__res[3];
  assign test_pe_comp__op_b[4] = test_opt_reg_file__res[4];
  assign test_pe_comp__op_b[5] = test_opt_reg_file__res[5];
  assign test_pe_comp__op_b[6] = test_opt_reg_file__res[6];
  assign test_pe_comp__op_b[7] = test_opt_reg_file__res[7];
  assign test_pe_comp__op_b[8] = test_opt_reg_file__res[8];
  assign test_pe_comp__op_b[9] = test_opt_reg_file__res[9];

endmodule //test_pe_unq1

module test_opt_reg_file (
  input [7:0] cfg_a,
  input [15:0] cfg_d,
  input  cfg_en,
  input  clk,
  input  clk_en,
  input [15:0] data_in,
  input  load,
  input [2:0] mode,
  output [15:0] reg_data,
  output [15:0] res,
  input  rst_n,
  input [15:0] val
);
  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89' (Module add_U11)
  wire [3:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B;
  wire [31:0] __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y;
  add_U11 __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89(
    .A(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A),
    .B(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B),
    .Y(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__Y)
  );

  //Wire declarations for instance '__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58' (Module and_U3)
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__A;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__B;
  wire [0:0] __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__Y;
  and_U3 __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58(
    .A(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__A),
    .B(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__B),
    .Y(__DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948' (Module reduce_or_U12)
  wire [2:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__Y;
  reduce_or_U12 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968' (Module reduce_or_U13)
  wire [1:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__Y;
  reduce_or_U13 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970' (Module not_U14)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970__Y;
  not_U14 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970__A),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964' (Module or_U6)
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__A;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__B;
  wire [0:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__Y;
  or_U6 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__B),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y)
  );

  //Wire declarations for instance '__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974' (Module rtMux_U10)
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B;
  wire  __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__S;
  wire [15:0] __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y;
  rtMux_U10 __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974(
    .A(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A),
    .B(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B),
    .S(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__S),
    .Y(__DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87' (Module eq_U15)
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A;
  wire [3:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__Y;
  eq_U15 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90' (Module eq_U16)
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A;
  wire [31:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__Y;
  eq_U16 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52' (Module eq_U17)
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A;
  wire [7:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__Y;
  eq_U17 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55' (Module eq_U18)
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__A;
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__Y;
  eq_U18 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57' (Module eq_U18)
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__A;
  wire [2:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__B;
  wire [0:0] __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__Y;
  eq_U18 __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57(
    .A(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__A),
    .B(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__B),
    .Y(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__Y)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__Y)
  );

  //Wire declarations for instance '__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51' (Module logic_and_U19)
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__A;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__B;
  wire [0:0] __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__Y;
  logic_and_U19 __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51(
    .A(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__A),
    .B(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__B),
    .Y(__DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__Y)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68' (Module lt_U20)
  wire [2:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__A;
  wire [31:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B;
  wire [0:0] __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__Y;
  lt_U20 __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68(
    .A(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__A),
    .B(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B),
    .Y(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__Y)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out)
  );

  //Wire declarations for instance '__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9' (Module corebit_const)
  wire  __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  corebit_const #(.value(0)) __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9(
    .out(__DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__Y)
  );

  //Wire declarations for instance '__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59' (Module or_U6)
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__A;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__B;
  wire [0:0] __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__Y;
  or_U6 __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59(
    .A(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__A),
    .B(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__B),
    .Y(__DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__Y)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__754' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__754__ARST;
  wire  __DOLLAR__procdff__DOLLAR__754__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__754__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__754__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__754(
    .ARST(__DOLLAR__procdff__DOLLAR__754__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__754__CLK),
    .D(__DOLLAR__procdff__DOLLAR__754__D),
    .Q(__DOLLAR__procdff__DOLLAR__754__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__755' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__755__ARST;
  wire  __DOLLAR__procdff__DOLLAR__755__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__755__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__755__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__755(
    .ARST(__DOLLAR__procdff__DOLLAR__755__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__755__CLK),
    .D(__DOLLAR__procdff__DOLLAR__755__D),
    .Q(__DOLLAR__procdff__DOLLAR__755__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__756' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__756__ARST;
  wire  __DOLLAR__procdff__DOLLAR__756__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__756__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__756__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__756(
    .ARST(__DOLLAR__procdff__DOLLAR__756__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__756__CLK),
    .D(__DOLLAR__procdff__DOLLAR__756__D),
    .Q(__DOLLAR__procdff__DOLLAR__756__Q)
  );

  //Wire declarations for instance '__DOLLAR__procdff__DOLLAR__757' (Module adff_U9)
  wire  __DOLLAR__procdff__DOLLAR__757__ARST;
  wire  __DOLLAR__procdff__DOLLAR__757__CLK;
  wire [15:0] __DOLLAR__procdff__DOLLAR__757__D;
  wire [15:0] __DOLLAR__procdff__DOLLAR__757__Q;
  adff_U9 #(.init(16'b0000000000000000)) __DOLLAR__procdff__DOLLAR__757(
    .ARST(__DOLLAR__procdff__DOLLAR__757__ARST),
    .CLK(__DOLLAR__procdff__DOLLAR__757__CLK),
    .D(__DOLLAR__procdff__DOLLAR__757__D),
    .Q(__DOLLAR__procdff__DOLLAR__757__Q)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__674' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__674__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__674__B;
  wire  __DOLLAR__procmux__DOLLAR__674__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__674__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__674(
    .A(__DOLLAR__procmux__DOLLAR__674__A),
    .B(__DOLLAR__procmux__DOLLAR__674__B),
    .S(__DOLLAR__procmux__DOLLAR__674__S),
    .Y(__DOLLAR__procmux__DOLLAR__674__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__677' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__677__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__677__B;
  wire  __DOLLAR__procmux__DOLLAR__677__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__677__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__677(
    .A(__DOLLAR__procmux__DOLLAR__677__A),
    .B(__DOLLAR__procmux__DOLLAR__677__B),
    .S(__DOLLAR__procmux__DOLLAR__677__S),
    .Y(__DOLLAR__procmux__DOLLAR__677__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__680' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__680__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__680__B;
  wire  __DOLLAR__procmux__DOLLAR__680__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__680__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__680(
    .A(__DOLLAR__procmux__DOLLAR__680__A),
    .B(__DOLLAR__procmux__DOLLAR__680__B),
    .S(__DOLLAR__procmux__DOLLAR__680__S),
    .Y(__DOLLAR__procmux__DOLLAR__680__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__684_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__684_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__684_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__684_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__684_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__684_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__684_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__685_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__685_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__685_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__685_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__685_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__685_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__685_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0' (Module eq_U17)
  wire [7:0] __DOLLAR__procmux__DOLLAR__686_CMP0__A;
  wire [7:0] __DOLLAR__procmux__DOLLAR__686_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__686_CMP0__Y;
  eq_U17 __DOLLAR__procmux__DOLLAR__686_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__686_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__686_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__686_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7(
    .out(__DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__689_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__689_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__689_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__689_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__689_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__689_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__689_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__689_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__690_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__690_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__690_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__690_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__690_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__690_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__690_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__690_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__691_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__691_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__691_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__691_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__691_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__691_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__691_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__691_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__692_CMP0' (Module eq_U5)
  wire [1:0] __DOLLAR__procmux__DOLLAR__692_CMP0__A;
  wire [1:0] __DOLLAR__procmux__DOLLAR__692_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__692_CMP0__Y;
  eq_U5 __DOLLAR__procmux__DOLLAR__692_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__692_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__692_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__692_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__693__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__693__B;
  wire  __DOLLAR__procmux__DOLLAR__693__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__693__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__693(
    .A(__DOLLAR__procmux__DOLLAR__693__A),
    .B(__DOLLAR__procmux__DOLLAR__693__B),
    .S(__DOLLAR__procmux__DOLLAR__693__S),
    .Y(__DOLLAR__procmux__DOLLAR__693__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9(
    .OUT(__DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__694_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__694_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__694_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__694_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__694_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__694_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__694_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__694_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__697_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__697_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__697_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__697_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__697_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__697_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__697_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__697_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__698_CMP0' (Module eq_U18)
  wire [2:0] __DOLLAR__procmux__DOLLAR__698_CMP0__A;
  wire [2:0] __DOLLAR__procmux__DOLLAR__698_CMP0__B;
  wire [0:0] __DOLLAR__procmux__DOLLAR__698_CMP0__Y;
  eq_U18 __DOLLAR__procmux__DOLLAR__698_CMP0(
    .A(__DOLLAR__procmux__DOLLAR__698_CMP0__A),
    .B(__DOLLAR__procmux__DOLLAR__698_CMP0__B),
    .Y(__DOLLAR__procmux__DOLLAR__698_CMP0__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0(
    .out(__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  corebit_const #(.value(1)) __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1(
    .out(__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2' (Module corebit_const)
  wire  __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  corebit_const #(.value(0)) __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2(
    .out(__DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__706' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__706__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__706__B;
  wire  __DOLLAR__procmux__DOLLAR__706__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__706__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__706(
    .A(__DOLLAR__procmux__DOLLAR__706__A),
    .B(__DOLLAR__procmux__DOLLAR__706__B),
    .S(__DOLLAR__procmux__DOLLAR__706__S),
    .Y(__DOLLAR__procmux__DOLLAR__706__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__709' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__709__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__709__B;
  wire  __DOLLAR__procmux__DOLLAR__709__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__709__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__709(
    .A(__DOLLAR__procmux__DOLLAR__709__A),
    .B(__DOLLAR__procmux__DOLLAR__709__B),
    .S(__DOLLAR__procmux__DOLLAR__709__S),
    .Y(__DOLLAR__procmux__DOLLAR__709__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__712__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__712__B;
  wire  __DOLLAR__procmux__DOLLAR__712__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__712__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__712(
    .A(__DOLLAR__procmux__DOLLAR__712__A),
    .B(__DOLLAR__procmux__DOLLAR__712__B),
    .S(__DOLLAR__procmux__DOLLAR__712__S),
    .Y(__DOLLAR__procmux__DOLLAR__712__Y)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9' (Module unknownBit)
  wire  __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  unknownBit __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9(
    .OUT(__DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT)
  );

  //Wire declarations for instance '__DOLLAR__procmux__DOLLAR__715' (Module rtMux_U10)
  wire [15:0] __DOLLAR__procmux__DOLLAR__715__A;
  wire [15:0] __DOLLAR__procmux__DOLLAR__715__B;
  wire  __DOLLAR__procmux__DOLLAR__715__S;
  wire [15:0] __DOLLAR__procmux__DOLLAR__715__Y;
  rtMux_U10 __DOLLAR__procmux__DOLLAR__715(
    .A(__DOLLAR__procmux__DOLLAR__715__A),
    .B(__DOLLAR__procmux__DOLLAR__715__B),
    .S(__DOLLAR__procmux__DOLLAR__715__S),
    .Y(__DOLLAR__procmux__DOLLAR__715__Y)
  );

  //Wire declarations for instance '__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69' (Module rtMux_U10)
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B;
  wire  __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__S;
  wire [15:0] __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y;
  rtMux_U10 __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69(
    .A(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A),
    .B(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B),
    .S(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__S),
    .Y(__DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y)
  );

  //All the connections
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__S = __DOLLAR__procmux__DOLLAR__684_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__S = __DOLLAR__procmux__DOLLAR__686_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__S = __DOLLAR__procmux__DOLLAR__689_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__S = __DOLLAR__procmux__DOLLAR__691_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__S = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__S = __DOLLAR__procmux__DOLLAR__698_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__S = __DOLLAR__procmux__DOLLAR__697_CMP0__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[10] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[11] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[12] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[13] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[14] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[15] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[16] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[17] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[18] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[19] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[20] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[21] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[22] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[23] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[24] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[25] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[26] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[27] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[28] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[29] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[30] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[31] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[8] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__A[9] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[3] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[4] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[5] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[6] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__B[7] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__B[1] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__B[2] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[0] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[10] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___bit_const_10__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[11] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___bit_const_11__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[12] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___bit_const_12__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[13] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___bit_const_13__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[14] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___bit_const_14__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[15] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___bit_const_15__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[16] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__16__RIGHT_BRACKET___bit_const_16__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[17] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__17__RIGHT_BRACKET___bit_const_17__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[18] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__18__RIGHT_BRACKET___bit_const_18__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[19] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__19__RIGHT_BRACKET___bit_const_19__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[1] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[20] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__20__RIGHT_BRACKET___bit_const_20__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[21] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__21__RIGHT_BRACKET___bit_const_21__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[22] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__22__RIGHT_BRACKET___bit_const_22__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[23] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__23__RIGHT_BRACKET___bit_const_23__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[24] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__24__RIGHT_BRACKET___bit_const_24__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[25] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__25__RIGHT_BRACKET___bit_const_25__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[26] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__26__RIGHT_BRACKET___bit_const_26__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[27] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__27__RIGHT_BRACKET___bit_const_27__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[28] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__28__RIGHT_BRACKET___bit_const_28__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[29] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__29__RIGHT_BRACKET___bit_const_29__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[2] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[30] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__30__RIGHT_BRACKET___bit_const_30__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[31] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__31__RIGHT_BRACKET___bit_const_31__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[3] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[4] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[5] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[6] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[7] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[8] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___bit_const_8__out;
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__B[9] = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___bit_const_9__out;
  assign __DOLLAR__procdff__DOLLAR__754__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__754__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__755__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__755__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__756__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__756__CLK = clk;
  assign __DOLLAR__procdff__DOLLAR__757__ARST = rst_n;
  assign __DOLLAR__procdff__DOLLAR__757__CLK = clk;
  assign __DOLLAR__procmux__DOLLAR__674__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__Y[0];
  assign __DOLLAR__procmux__DOLLAR__677__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__Y[0];
  assign __DOLLAR__procmux__DOLLAR__680__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__Y[0];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__684_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__685_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[3] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___bit_const_3__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[4] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___bit_const_4__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[5] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___bit_const_5__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[6] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___bit_const_6__out;
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__B[7] = __DOLLAR__procmux__DOLLAR__686_CMP0__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___bit_const_7__out;
  assign __DOLLAR__procmux__DOLLAR__689_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__689_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__689_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__690_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__690_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__690_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__691_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__691_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__691_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__692_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__692_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__692_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__693__S = __DOLLAR__procmux__DOLLAR__694_CMP0__Y[0];
  assign __DOLLAR__procmux__DOLLAR__693__A[0] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[10] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[11] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[12] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[13] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[14] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[15] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[1] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[2] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[3] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[4] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[5] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[6] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[7] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[8] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  assign __DOLLAR__procmux__DOLLAR__693__A[9] = __DOLLAR__procmux__DOLLAR__693__DOT__A__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__694_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__697_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__B[0] = __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___bit_const_0__out;
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__B[1] = __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___bit_const_1__out;
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__B[2] = __DOLLAR__procmux__DOLLAR__698_CMP0__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___bit_const_2__out;
  assign __DOLLAR__procmux__DOLLAR__706__S = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__Y[0];
  assign __DOLLAR__procmux__DOLLAR__709__S = load;
  assign __DOLLAR__procmux__DOLLAR__712__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__Y[0];
  assign __DOLLAR__procmux__DOLLAR__712__B[0] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__0__RIGHT_BRACKET___unknown_value_0__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[10] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__10__RIGHT_BRACKET___unknown_value_10__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[11] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__11__RIGHT_BRACKET___unknown_value_11__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[12] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__12__RIGHT_BRACKET___unknown_value_12__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[13] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__13__RIGHT_BRACKET___unknown_value_13__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[14] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__14__RIGHT_BRACKET___unknown_value_14__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[15] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__15__RIGHT_BRACKET___unknown_value_15__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[1] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__1__RIGHT_BRACKET___unknown_value_1__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[2] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__2__RIGHT_BRACKET___unknown_value_2__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[3] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__3__RIGHT_BRACKET___unknown_value_3__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[4] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__4__RIGHT_BRACKET___unknown_value_4__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[5] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__5__RIGHT_BRACKET___unknown_value_5__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[6] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__6__RIGHT_BRACKET___unknown_value_6__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[7] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__7__RIGHT_BRACKET___unknown_value_7__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[8] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__8__RIGHT_BRACKET___unknown_value_8__OUT;
  assign __DOLLAR__procmux__DOLLAR__712__B[9] = __DOLLAR__procmux__DOLLAR__712__DOT__B__LEFT_BRACKET__9__RIGHT_BRACKET___unknown_value_9__OUT;
  assign __DOLLAR__procmux__DOLLAR__715__S = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__S = __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__A[0] = cfg_en;
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__A[0] = cfg_en;
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__B[0] = clk_en;
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__A[0] = load;
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__75__Y[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__82__Y[9];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A[0] = cfg_a[0];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A[1] = cfg_a[1];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A[2] = cfg_a[2];
  assign __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[0] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[1] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[10] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[10];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[11] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[11];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[12] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[12];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[13] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[13];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[14] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[14];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[15] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[15];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[16] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[16];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[17] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[17];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[18] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[18];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[19] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[19];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[2] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[20] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[20];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[21] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[21];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[22] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[22];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[23] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[23];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[24] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[24];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[25] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[25];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[26] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[26];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[27] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[27];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[28] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[28];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[29] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[29];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[3] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[30] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[30];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[31] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[31];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[4] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[5] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[6] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[7] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[8] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[8];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__B[9] = __DOLLAR__add__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__89__Y[9];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__53__Y[0];
  assign __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__A[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__B[0] = __DOLLAR__and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__58__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__A[0] = __DOLLAR__procmux__DOLLAR__684_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__A[1] = __DOLLAR__procmux__DOLLAR__685_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__A[2] = __DOLLAR__procmux__DOLLAR__686_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__950__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__948__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__A[0] = __DOLLAR__procmux__DOLLAR__697_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__A[1] = __DOLLAR__procmux__DOLLAR__698_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__101__COLON__execute__DOLLAR__970__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__100__COLON__execute__DOLLAR__968__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__A[0] = __DOLLAR__procmux__DOLLAR__685_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__956__B[0] = __DOLLAR__procmux__DOLLAR__684_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__A[0] = __DOLLAR__procmux__DOLLAR__690_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__35__COLON__or_generator__DOLLAR__964__B[0] = __DOLLAR__procmux__DOLLAR__689_CMP0__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[0] = __DOLLAR__procdff__DOLLAR__755__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[1] = __DOLLAR__procdff__DOLLAR__755__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[10] = __DOLLAR__procdff__DOLLAR__755__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[11] = __DOLLAR__procdff__DOLLAR__755__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[12] = __DOLLAR__procdff__DOLLAR__755__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[13] = __DOLLAR__procdff__DOLLAR__755__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[14] = __DOLLAR__procdff__DOLLAR__755__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[15] = __DOLLAR__procdff__DOLLAR__755__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[2] = __DOLLAR__procdff__DOLLAR__755__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[3] = __DOLLAR__procdff__DOLLAR__755__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[4] = __DOLLAR__procdff__DOLLAR__755__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[5] = __DOLLAR__procdff__DOLLAR__755__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[6] = __DOLLAR__procdff__DOLLAR__755__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[7] = __DOLLAR__procdff__DOLLAR__755__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[8] = __DOLLAR__procdff__DOLLAR__755__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__A[9] = __DOLLAR__procdff__DOLLAR__755__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[0] = __DOLLAR__procdff__DOLLAR__754__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[1] = __DOLLAR__procdff__DOLLAR__754__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[10] = __DOLLAR__procdff__DOLLAR__754__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[11] = __DOLLAR__procdff__DOLLAR__754__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[12] = __DOLLAR__procdff__DOLLAR__754__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[13] = __DOLLAR__procdff__DOLLAR__754__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[14] = __DOLLAR__procdff__DOLLAR__754__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[15] = __DOLLAR__procdff__DOLLAR__754__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[2] = __DOLLAR__procdff__DOLLAR__754__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[3] = __DOLLAR__procdff__DOLLAR__754__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[4] = __DOLLAR__procdff__DOLLAR__754__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[5] = __DOLLAR__procdff__DOLLAR__754__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[6] = __DOLLAR__procdff__DOLLAR__754__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[7] = __DOLLAR__procdff__DOLLAR__754__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[8] = __DOLLAR__procdff__DOLLAR__754__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__B[9] = __DOLLAR__procdff__DOLLAR__754__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__952__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[0] = __DOLLAR__procdff__DOLLAR__757__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[1] = __DOLLAR__procdff__DOLLAR__757__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[10] = __DOLLAR__procdff__DOLLAR__757__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[11] = __DOLLAR__procdff__DOLLAR__757__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[12] = __DOLLAR__procdff__DOLLAR__757__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[13] = __DOLLAR__procdff__DOLLAR__757__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[14] = __DOLLAR__procdff__DOLLAR__757__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[15] = __DOLLAR__procdff__DOLLAR__757__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[2] = __DOLLAR__procdff__DOLLAR__757__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[3] = __DOLLAR__procdff__DOLLAR__757__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[4] = __DOLLAR__procdff__DOLLAR__757__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[5] = __DOLLAR__procdff__DOLLAR__757__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[6] = __DOLLAR__procdff__DOLLAR__757__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[7] = __DOLLAR__procdff__DOLLAR__757__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[8] = __DOLLAR__procdff__DOLLAR__757__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__A[9] = __DOLLAR__procdff__DOLLAR__757__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[0] = __DOLLAR__procdff__DOLLAR__756__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[1] = __DOLLAR__procdff__DOLLAR__756__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[10] = __DOLLAR__procdff__DOLLAR__756__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[11] = __DOLLAR__procdff__DOLLAR__756__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[12] = __DOLLAR__procdff__DOLLAR__756__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[13] = __DOLLAR__procdff__DOLLAR__756__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[14] = __DOLLAR__procdff__DOLLAR__756__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[15] = __DOLLAR__procdff__DOLLAR__756__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[2] = __DOLLAR__procdff__DOLLAR__756__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[3] = __DOLLAR__procdff__DOLLAR__756__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[4] = __DOLLAR__procdff__DOLLAR__756__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[5] = __DOLLAR__procdff__DOLLAR__756__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[6] = __DOLLAR__procdff__DOLLAR__756__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[7] = __DOLLAR__procdff__DOLLAR__756__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[8] = __DOLLAR__procdff__DOLLAR__756__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__B[9] = __DOLLAR__procdff__DOLLAR__756__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__954__Y[9];
  assign reg_data[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[0];
  assign reg_data[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[1];
  assign reg_data[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[10];
  assign reg_data[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[11];
  assign reg_data[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[12];
  assign reg_data[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[13];
  assign reg_data[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[14];
  assign reg_data[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[15];
  assign reg_data[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[2];
  assign reg_data[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[3];
  assign reg_data[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[4];
  assign reg_data[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[5];
  assign reg_data[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[6];
  assign reg_data[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[7];
  assign reg_data[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[8];
  assign reg_data[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__958__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[0] = __DOLLAR__procdff__DOLLAR__755__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[1] = __DOLLAR__procdff__DOLLAR__755__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[10] = __DOLLAR__procdff__DOLLAR__755__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[11] = __DOLLAR__procdff__DOLLAR__755__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[12] = __DOLLAR__procdff__DOLLAR__755__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[13] = __DOLLAR__procdff__DOLLAR__755__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[14] = __DOLLAR__procdff__DOLLAR__755__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[15] = __DOLLAR__procdff__DOLLAR__755__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[2] = __DOLLAR__procdff__DOLLAR__755__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[3] = __DOLLAR__procdff__DOLLAR__755__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[4] = __DOLLAR__procdff__DOLLAR__755__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[5] = __DOLLAR__procdff__DOLLAR__755__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[6] = __DOLLAR__procdff__DOLLAR__755__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[7] = __DOLLAR__procdff__DOLLAR__755__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[8] = __DOLLAR__procdff__DOLLAR__755__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__A[9] = __DOLLAR__procdff__DOLLAR__755__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[0] = __DOLLAR__procdff__DOLLAR__754__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[1] = __DOLLAR__procdff__DOLLAR__754__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[10] = __DOLLAR__procdff__DOLLAR__754__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[11] = __DOLLAR__procdff__DOLLAR__754__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[12] = __DOLLAR__procdff__DOLLAR__754__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[13] = __DOLLAR__procdff__DOLLAR__754__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[14] = __DOLLAR__procdff__DOLLAR__754__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[15] = __DOLLAR__procdff__DOLLAR__754__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[2] = __DOLLAR__procdff__DOLLAR__754__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[3] = __DOLLAR__procdff__DOLLAR__754__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[4] = __DOLLAR__procdff__DOLLAR__754__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[5] = __DOLLAR__procdff__DOLLAR__754__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[6] = __DOLLAR__procdff__DOLLAR__754__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[7] = __DOLLAR__procdff__DOLLAR__754__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[8] = __DOLLAR__procdff__DOLLAR__754__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__B[9] = __DOLLAR__procdff__DOLLAR__754__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__960__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[0] = __DOLLAR__procdff__DOLLAR__757__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[1] = __DOLLAR__procdff__DOLLAR__757__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[10] = __DOLLAR__procdff__DOLLAR__757__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[11] = __DOLLAR__procdff__DOLLAR__757__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[12] = __DOLLAR__procdff__DOLLAR__757__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[13] = __DOLLAR__procdff__DOLLAR__757__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[14] = __DOLLAR__procdff__DOLLAR__757__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[15] = __DOLLAR__procdff__DOLLAR__757__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[2] = __DOLLAR__procdff__DOLLAR__757__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[3] = __DOLLAR__procdff__DOLLAR__757__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[4] = __DOLLAR__procdff__DOLLAR__757__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[5] = __DOLLAR__procdff__DOLLAR__757__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[6] = __DOLLAR__procdff__DOLLAR__757__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[7] = __DOLLAR__procdff__DOLLAR__757__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[8] = __DOLLAR__procdff__DOLLAR__757__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__A[9] = __DOLLAR__procdff__DOLLAR__757__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[0] = __DOLLAR__procdff__DOLLAR__756__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[1] = __DOLLAR__procdff__DOLLAR__756__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[10] = __DOLLAR__procdff__DOLLAR__756__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[11] = __DOLLAR__procdff__DOLLAR__756__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[12] = __DOLLAR__procdff__DOLLAR__756__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[13] = __DOLLAR__procdff__DOLLAR__756__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[14] = __DOLLAR__procdff__DOLLAR__756__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[15] = __DOLLAR__procdff__DOLLAR__756__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[2] = __DOLLAR__procdff__DOLLAR__756__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[3] = __DOLLAR__procdff__DOLLAR__756__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[4] = __DOLLAR__procdff__DOLLAR__756__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[5] = __DOLLAR__procdff__DOLLAR__756__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[6] = __DOLLAR__procdff__DOLLAR__756__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[7] = __DOLLAR__procdff__DOLLAR__756__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[8] = __DOLLAR__procdff__DOLLAR__756__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__B[9] = __DOLLAR__procdff__DOLLAR__756__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__962__Y[9];
  assign __DOLLAR__procmux__DOLLAR__693__B[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[0];
  assign __DOLLAR__procmux__DOLLAR__693__B[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[1];
  assign __DOLLAR__procmux__DOLLAR__693__B[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[10];
  assign __DOLLAR__procmux__DOLLAR__693__B[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[11];
  assign __DOLLAR__procmux__DOLLAR__693__B[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[12];
  assign __DOLLAR__procmux__DOLLAR__693__B[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[13];
  assign __DOLLAR__procmux__DOLLAR__693__B[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[14];
  assign __DOLLAR__procmux__DOLLAR__693__B[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[15];
  assign __DOLLAR__procmux__DOLLAR__693__B[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[2];
  assign __DOLLAR__procmux__DOLLAR__693__B[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[3];
  assign __DOLLAR__procmux__DOLLAR__693__B[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[4];
  assign __DOLLAR__procmux__DOLLAR__693__B[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[5];
  assign __DOLLAR__procmux__DOLLAR__693__B[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[6];
  assign __DOLLAR__procmux__DOLLAR__693__B[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[7];
  assign __DOLLAR__procmux__DOLLAR__693__B[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[8];
  assign __DOLLAR__procmux__DOLLAR__693__B[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__966__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[0] = __DOLLAR__procdff__DOLLAR__757__Q[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[1] = __DOLLAR__procdff__DOLLAR__757__Q[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[10] = __DOLLAR__procdff__DOLLAR__757__Q[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[11] = __DOLLAR__procdff__DOLLAR__757__Q[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[12] = __DOLLAR__procdff__DOLLAR__757__Q[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[13] = __DOLLAR__procdff__DOLLAR__757__Q[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[14] = __DOLLAR__procdff__DOLLAR__757__Q[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[15] = __DOLLAR__procdff__DOLLAR__757__Q[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[2] = __DOLLAR__procdff__DOLLAR__757__Q[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[3] = __DOLLAR__procdff__DOLLAR__757__Q[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[4] = __DOLLAR__procdff__DOLLAR__757__Q[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[5] = __DOLLAR__procdff__DOLLAR__757__Q[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[6] = __DOLLAR__procdff__DOLLAR__757__Q[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[7] = __DOLLAR__procdff__DOLLAR__757__Q[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[8] = __DOLLAR__procdff__DOLLAR__757__Q[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__A[9] = __DOLLAR__procdff__DOLLAR__757__Q[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[0] = data_in[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[1] = data_in[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[10] = data_in[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[11] = data_in[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[12] = data_in[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[13] = data_in[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[14] = data_in[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[15] = data_in[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[2] = data_in[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[3] = data_in[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[4] = data_in[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[5] = data_in[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[6] = data_in[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[7] = data_in[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[8] = data_in[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__B[9] = data_in[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__A[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__972__Y[9];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[0] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[0];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[1] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[1];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[10] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[10];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[11] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[11];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[12] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[12];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[13] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[13];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[14] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[14];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[15] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[15];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[2] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[2];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[3] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[3];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[4] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[4];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[5] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[5];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[6] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[6];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[7] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[7];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[8] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[8];
  assign __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__B[9] = __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__Y[9];
  assign res[0] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[0];
  assign res[1] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[1];
  assign res[10] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[10];
  assign res[11] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[11];
  assign res[12] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[12];
  assign res[13] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[13];
  assign res[14] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[14];
  assign res[15] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[15];
  assign res[2] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[2];
  assign res[3] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[3];
  assign res[4] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[4];
  assign res[5] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[5];
  assign res[6] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[6];
  assign res[7] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[7];
  assign res[8] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[8];
  assign res[9] = __DOLLAR__auto__DOLLAR__pmuxtree__DOT__cc__COLON__65__COLON__recursive_mux_generator__DOLLAR__974__Y[9];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__73__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__76__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__80__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__83__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A[0] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A[1] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A[2] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__A[3] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__87__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__90__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__A[7] = cfg_a[7];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__51__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__74__DOLLAR__50__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[0] = cfg_a[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[1] = cfg_a[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[2] = cfg_a[2];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[3] = cfg_a[3];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[4] = cfg_a[4];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[5] = cfg_a[5];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[6] = cfg_a[6];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__52__A[7] = cfg_a[7];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__A[2] = mode[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__B[0] = __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__55__Y[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__A[0] = mode[0];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__A[1] = mode[1];
  assign __DOLLAR__eq__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__57__A[2] = mode[2];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__77__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__74__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__84__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__81__Y[0];
  assign __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__91__A[0] = __DOLLAR__logic_and__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__104__DOLLAR__88__Y[0];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__A[0] = data_in[0];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__A[1] = data_in[1];
  assign __DOLLAR__lt__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__117__DOLLAR__68__A[2] = data_in[2];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__84__DOLLAR__54__Y[0];
  assign __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__86__DOLLAR__59__A[0] = __DOLLAR__or__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__85__DOLLAR__56__Y[0];
  assign __DOLLAR__procdff__DOLLAR__754__D[0] = __DOLLAR__procmux__DOLLAR__674__Y[0];
  assign __DOLLAR__procdff__DOLLAR__754__D[1] = __DOLLAR__procmux__DOLLAR__674__Y[1];
  assign __DOLLAR__procdff__DOLLAR__754__D[10] = __DOLLAR__procmux__DOLLAR__674__Y[10];
  assign __DOLLAR__procdff__DOLLAR__754__D[11] = __DOLLAR__procmux__DOLLAR__674__Y[11];
  assign __DOLLAR__procdff__DOLLAR__754__D[12] = __DOLLAR__procmux__DOLLAR__674__Y[12];
  assign __DOLLAR__procdff__DOLLAR__754__D[13] = __DOLLAR__procmux__DOLLAR__674__Y[13];
  assign __DOLLAR__procdff__DOLLAR__754__D[14] = __DOLLAR__procmux__DOLLAR__674__Y[14];
  assign __DOLLAR__procdff__DOLLAR__754__D[15] = __DOLLAR__procmux__DOLLAR__674__Y[15];
  assign __DOLLAR__procdff__DOLLAR__754__D[2] = __DOLLAR__procmux__DOLLAR__674__Y[2];
  assign __DOLLAR__procdff__DOLLAR__754__D[3] = __DOLLAR__procmux__DOLLAR__674__Y[3];
  assign __DOLLAR__procdff__DOLLAR__754__D[4] = __DOLLAR__procmux__DOLLAR__674__Y[4];
  assign __DOLLAR__procdff__DOLLAR__754__D[5] = __DOLLAR__procmux__DOLLAR__674__Y[5];
  assign __DOLLAR__procdff__DOLLAR__754__D[6] = __DOLLAR__procmux__DOLLAR__674__Y[6];
  assign __DOLLAR__procdff__DOLLAR__754__D[7] = __DOLLAR__procmux__DOLLAR__674__Y[7];
  assign __DOLLAR__procdff__DOLLAR__754__D[8] = __DOLLAR__procmux__DOLLAR__674__Y[8];
  assign __DOLLAR__procdff__DOLLAR__754__D[9] = __DOLLAR__procmux__DOLLAR__674__Y[9];
  assign __DOLLAR__procmux__DOLLAR__674__A[0] = __DOLLAR__procdff__DOLLAR__754__Q[0];
  assign __DOLLAR__procmux__DOLLAR__674__A[1] = __DOLLAR__procdff__DOLLAR__754__Q[1];
  assign __DOLLAR__procmux__DOLLAR__674__A[10] = __DOLLAR__procdff__DOLLAR__754__Q[10];
  assign __DOLLAR__procmux__DOLLAR__674__A[11] = __DOLLAR__procdff__DOLLAR__754__Q[11];
  assign __DOLLAR__procmux__DOLLAR__674__A[12] = __DOLLAR__procdff__DOLLAR__754__Q[12];
  assign __DOLLAR__procmux__DOLLAR__674__A[13] = __DOLLAR__procdff__DOLLAR__754__Q[13];
  assign __DOLLAR__procmux__DOLLAR__674__A[14] = __DOLLAR__procdff__DOLLAR__754__Q[14];
  assign __DOLLAR__procmux__DOLLAR__674__A[15] = __DOLLAR__procdff__DOLLAR__754__Q[15];
  assign __DOLLAR__procmux__DOLLAR__674__A[2] = __DOLLAR__procdff__DOLLAR__754__Q[2];
  assign __DOLLAR__procmux__DOLLAR__674__A[3] = __DOLLAR__procdff__DOLLAR__754__Q[3];
  assign __DOLLAR__procmux__DOLLAR__674__A[4] = __DOLLAR__procdff__DOLLAR__754__Q[4];
  assign __DOLLAR__procmux__DOLLAR__674__A[5] = __DOLLAR__procdff__DOLLAR__754__Q[5];
  assign __DOLLAR__procmux__DOLLAR__674__A[6] = __DOLLAR__procdff__DOLLAR__754__Q[6];
  assign __DOLLAR__procmux__DOLLAR__674__A[7] = __DOLLAR__procdff__DOLLAR__754__Q[7];
  assign __DOLLAR__procmux__DOLLAR__674__A[8] = __DOLLAR__procdff__DOLLAR__754__Q[8];
  assign __DOLLAR__procmux__DOLLAR__674__A[9] = __DOLLAR__procdff__DOLLAR__754__Q[9];
  assign __DOLLAR__procdff__DOLLAR__755__D[0] = __DOLLAR__procmux__DOLLAR__677__Y[0];
  assign __DOLLAR__procdff__DOLLAR__755__D[1] = __DOLLAR__procmux__DOLLAR__677__Y[1];
  assign __DOLLAR__procdff__DOLLAR__755__D[10] = __DOLLAR__procmux__DOLLAR__677__Y[10];
  assign __DOLLAR__procdff__DOLLAR__755__D[11] = __DOLLAR__procmux__DOLLAR__677__Y[11];
  assign __DOLLAR__procdff__DOLLAR__755__D[12] = __DOLLAR__procmux__DOLLAR__677__Y[12];
  assign __DOLLAR__procdff__DOLLAR__755__D[13] = __DOLLAR__procmux__DOLLAR__677__Y[13];
  assign __DOLLAR__procdff__DOLLAR__755__D[14] = __DOLLAR__procmux__DOLLAR__677__Y[14];
  assign __DOLLAR__procdff__DOLLAR__755__D[15] = __DOLLAR__procmux__DOLLAR__677__Y[15];
  assign __DOLLAR__procdff__DOLLAR__755__D[2] = __DOLLAR__procmux__DOLLAR__677__Y[2];
  assign __DOLLAR__procdff__DOLLAR__755__D[3] = __DOLLAR__procmux__DOLLAR__677__Y[3];
  assign __DOLLAR__procdff__DOLLAR__755__D[4] = __DOLLAR__procmux__DOLLAR__677__Y[4];
  assign __DOLLAR__procdff__DOLLAR__755__D[5] = __DOLLAR__procmux__DOLLAR__677__Y[5];
  assign __DOLLAR__procdff__DOLLAR__755__D[6] = __DOLLAR__procmux__DOLLAR__677__Y[6];
  assign __DOLLAR__procdff__DOLLAR__755__D[7] = __DOLLAR__procmux__DOLLAR__677__Y[7];
  assign __DOLLAR__procdff__DOLLAR__755__D[8] = __DOLLAR__procmux__DOLLAR__677__Y[8];
  assign __DOLLAR__procdff__DOLLAR__755__D[9] = __DOLLAR__procmux__DOLLAR__677__Y[9];
  assign __DOLLAR__procmux__DOLLAR__677__A[0] = __DOLLAR__procdff__DOLLAR__755__Q[0];
  assign __DOLLAR__procmux__DOLLAR__677__A[1] = __DOLLAR__procdff__DOLLAR__755__Q[1];
  assign __DOLLAR__procmux__DOLLAR__677__A[10] = __DOLLAR__procdff__DOLLAR__755__Q[10];
  assign __DOLLAR__procmux__DOLLAR__677__A[11] = __DOLLAR__procdff__DOLLAR__755__Q[11];
  assign __DOLLAR__procmux__DOLLAR__677__A[12] = __DOLLAR__procdff__DOLLAR__755__Q[12];
  assign __DOLLAR__procmux__DOLLAR__677__A[13] = __DOLLAR__procdff__DOLLAR__755__Q[13];
  assign __DOLLAR__procmux__DOLLAR__677__A[14] = __DOLLAR__procdff__DOLLAR__755__Q[14];
  assign __DOLLAR__procmux__DOLLAR__677__A[15] = __DOLLAR__procdff__DOLLAR__755__Q[15];
  assign __DOLLAR__procmux__DOLLAR__677__A[2] = __DOLLAR__procdff__DOLLAR__755__Q[2];
  assign __DOLLAR__procmux__DOLLAR__677__A[3] = __DOLLAR__procdff__DOLLAR__755__Q[3];
  assign __DOLLAR__procmux__DOLLAR__677__A[4] = __DOLLAR__procdff__DOLLAR__755__Q[4];
  assign __DOLLAR__procmux__DOLLAR__677__A[5] = __DOLLAR__procdff__DOLLAR__755__Q[5];
  assign __DOLLAR__procmux__DOLLAR__677__A[6] = __DOLLAR__procdff__DOLLAR__755__Q[6];
  assign __DOLLAR__procmux__DOLLAR__677__A[7] = __DOLLAR__procdff__DOLLAR__755__Q[7];
  assign __DOLLAR__procmux__DOLLAR__677__A[8] = __DOLLAR__procdff__DOLLAR__755__Q[8];
  assign __DOLLAR__procmux__DOLLAR__677__A[9] = __DOLLAR__procdff__DOLLAR__755__Q[9];
  assign __DOLLAR__procdff__DOLLAR__756__D[0] = __DOLLAR__procmux__DOLLAR__680__Y[0];
  assign __DOLLAR__procdff__DOLLAR__756__D[1] = __DOLLAR__procmux__DOLLAR__680__Y[1];
  assign __DOLLAR__procdff__DOLLAR__756__D[10] = __DOLLAR__procmux__DOLLAR__680__Y[10];
  assign __DOLLAR__procdff__DOLLAR__756__D[11] = __DOLLAR__procmux__DOLLAR__680__Y[11];
  assign __DOLLAR__procdff__DOLLAR__756__D[12] = __DOLLAR__procmux__DOLLAR__680__Y[12];
  assign __DOLLAR__procdff__DOLLAR__756__D[13] = __DOLLAR__procmux__DOLLAR__680__Y[13];
  assign __DOLLAR__procdff__DOLLAR__756__D[14] = __DOLLAR__procmux__DOLLAR__680__Y[14];
  assign __DOLLAR__procdff__DOLLAR__756__D[15] = __DOLLAR__procmux__DOLLAR__680__Y[15];
  assign __DOLLAR__procdff__DOLLAR__756__D[2] = __DOLLAR__procmux__DOLLAR__680__Y[2];
  assign __DOLLAR__procdff__DOLLAR__756__D[3] = __DOLLAR__procmux__DOLLAR__680__Y[3];
  assign __DOLLAR__procdff__DOLLAR__756__D[4] = __DOLLAR__procmux__DOLLAR__680__Y[4];
  assign __DOLLAR__procdff__DOLLAR__756__D[5] = __DOLLAR__procmux__DOLLAR__680__Y[5];
  assign __DOLLAR__procdff__DOLLAR__756__D[6] = __DOLLAR__procmux__DOLLAR__680__Y[6];
  assign __DOLLAR__procdff__DOLLAR__756__D[7] = __DOLLAR__procmux__DOLLAR__680__Y[7];
  assign __DOLLAR__procdff__DOLLAR__756__D[8] = __DOLLAR__procmux__DOLLAR__680__Y[8];
  assign __DOLLAR__procdff__DOLLAR__756__D[9] = __DOLLAR__procmux__DOLLAR__680__Y[9];
  assign __DOLLAR__procmux__DOLLAR__680__A[0] = __DOLLAR__procdff__DOLLAR__756__Q[0];
  assign __DOLLAR__procmux__DOLLAR__680__A[1] = __DOLLAR__procdff__DOLLAR__756__Q[1];
  assign __DOLLAR__procmux__DOLLAR__680__A[10] = __DOLLAR__procdff__DOLLAR__756__Q[10];
  assign __DOLLAR__procmux__DOLLAR__680__A[11] = __DOLLAR__procdff__DOLLAR__756__Q[11];
  assign __DOLLAR__procmux__DOLLAR__680__A[12] = __DOLLAR__procdff__DOLLAR__756__Q[12];
  assign __DOLLAR__procmux__DOLLAR__680__A[13] = __DOLLAR__procdff__DOLLAR__756__Q[13];
  assign __DOLLAR__procmux__DOLLAR__680__A[14] = __DOLLAR__procdff__DOLLAR__756__Q[14];
  assign __DOLLAR__procmux__DOLLAR__680__A[15] = __DOLLAR__procdff__DOLLAR__756__Q[15];
  assign __DOLLAR__procmux__DOLLAR__680__A[2] = __DOLLAR__procdff__DOLLAR__756__Q[2];
  assign __DOLLAR__procmux__DOLLAR__680__A[3] = __DOLLAR__procdff__DOLLAR__756__Q[3];
  assign __DOLLAR__procmux__DOLLAR__680__A[4] = __DOLLAR__procdff__DOLLAR__756__Q[4];
  assign __DOLLAR__procmux__DOLLAR__680__A[5] = __DOLLAR__procdff__DOLLAR__756__Q[5];
  assign __DOLLAR__procmux__DOLLAR__680__A[6] = __DOLLAR__procdff__DOLLAR__756__Q[6];
  assign __DOLLAR__procmux__DOLLAR__680__A[7] = __DOLLAR__procdff__DOLLAR__756__Q[7];
  assign __DOLLAR__procmux__DOLLAR__680__A[8] = __DOLLAR__procdff__DOLLAR__756__Q[8];
  assign __DOLLAR__procmux__DOLLAR__680__A[9] = __DOLLAR__procdff__DOLLAR__756__Q[9];
  assign __DOLLAR__procdff__DOLLAR__757__D[0] = __DOLLAR__procmux__DOLLAR__706__Y[0];
  assign __DOLLAR__procdff__DOLLAR__757__D[1] = __DOLLAR__procmux__DOLLAR__706__Y[1];
  assign __DOLLAR__procdff__DOLLAR__757__D[10] = __DOLLAR__procmux__DOLLAR__706__Y[10];
  assign __DOLLAR__procdff__DOLLAR__757__D[11] = __DOLLAR__procmux__DOLLAR__706__Y[11];
  assign __DOLLAR__procdff__DOLLAR__757__D[12] = __DOLLAR__procmux__DOLLAR__706__Y[12];
  assign __DOLLAR__procdff__DOLLAR__757__D[13] = __DOLLAR__procmux__DOLLAR__706__Y[13];
  assign __DOLLAR__procdff__DOLLAR__757__D[14] = __DOLLAR__procmux__DOLLAR__706__Y[14];
  assign __DOLLAR__procdff__DOLLAR__757__D[15] = __DOLLAR__procmux__DOLLAR__706__Y[15];
  assign __DOLLAR__procdff__DOLLAR__757__D[2] = __DOLLAR__procmux__DOLLAR__706__Y[2];
  assign __DOLLAR__procdff__DOLLAR__757__D[3] = __DOLLAR__procmux__DOLLAR__706__Y[3];
  assign __DOLLAR__procdff__DOLLAR__757__D[4] = __DOLLAR__procmux__DOLLAR__706__Y[4];
  assign __DOLLAR__procdff__DOLLAR__757__D[5] = __DOLLAR__procmux__DOLLAR__706__Y[5];
  assign __DOLLAR__procdff__DOLLAR__757__D[6] = __DOLLAR__procmux__DOLLAR__706__Y[6];
  assign __DOLLAR__procdff__DOLLAR__757__D[7] = __DOLLAR__procmux__DOLLAR__706__Y[7];
  assign __DOLLAR__procdff__DOLLAR__757__D[8] = __DOLLAR__procmux__DOLLAR__706__Y[8];
  assign __DOLLAR__procdff__DOLLAR__757__D[9] = __DOLLAR__procmux__DOLLAR__706__Y[9];
  assign __DOLLAR__procmux__DOLLAR__706__A[0] = __DOLLAR__procdff__DOLLAR__757__Q[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[0] = __DOLLAR__procdff__DOLLAR__757__Q[0];
  assign __DOLLAR__procmux__DOLLAR__706__A[1] = __DOLLAR__procdff__DOLLAR__757__Q[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[1] = __DOLLAR__procdff__DOLLAR__757__Q[1];
  assign __DOLLAR__procmux__DOLLAR__706__A[10] = __DOLLAR__procdff__DOLLAR__757__Q[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[10] = __DOLLAR__procdff__DOLLAR__757__Q[10];
  assign __DOLLAR__procmux__DOLLAR__706__A[11] = __DOLLAR__procdff__DOLLAR__757__Q[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[11] = __DOLLAR__procdff__DOLLAR__757__Q[11];
  assign __DOLLAR__procmux__DOLLAR__706__A[12] = __DOLLAR__procdff__DOLLAR__757__Q[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[12] = __DOLLAR__procdff__DOLLAR__757__Q[12];
  assign __DOLLAR__procmux__DOLLAR__706__A[13] = __DOLLAR__procdff__DOLLAR__757__Q[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[13] = __DOLLAR__procdff__DOLLAR__757__Q[13];
  assign __DOLLAR__procmux__DOLLAR__706__A[14] = __DOLLAR__procdff__DOLLAR__757__Q[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[14] = __DOLLAR__procdff__DOLLAR__757__Q[14];
  assign __DOLLAR__procmux__DOLLAR__706__A[15] = __DOLLAR__procdff__DOLLAR__757__Q[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[15] = __DOLLAR__procdff__DOLLAR__757__Q[15];
  assign __DOLLAR__procmux__DOLLAR__706__A[2] = __DOLLAR__procdff__DOLLAR__757__Q[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[2] = __DOLLAR__procdff__DOLLAR__757__Q[2];
  assign __DOLLAR__procmux__DOLLAR__706__A[3] = __DOLLAR__procdff__DOLLAR__757__Q[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[3] = __DOLLAR__procdff__DOLLAR__757__Q[3];
  assign __DOLLAR__procmux__DOLLAR__706__A[4] = __DOLLAR__procdff__DOLLAR__757__Q[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[4] = __DOLLAR__procdff__DOLLAR__757__Q[4];
  assign __DOLLAR__procmux__DOLLAR__706__A[5] = __DOLLAR__procdff__DOLLAR__757__Q[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[5] = __DOLLAR__procdff__DOLLAR__757__Q[5];
  assign __DOLLAR__procmux__DOLLAR__706__A[6] = __DOLLAR__procdff__DOLLAR__757__Q[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[6] = __DOLLAR__procdff__DOLLAR__757__Q[6];
  assign __DOLLAR__procmux__DOLLAR__706__A[7] = __DOLLAR__procdff__DOLLAR__757__Q[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[7] = __DOLLAR__procdff__DOLLAR__757__Q[7];
  assign __DOLLAR__procmux__DOLLAR__706__A[8] = __DOLLAR__procdff__DOLLAR__757__Q[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[8] = __DOLLAR__procdff__DOLLAR__757__Q[8];
  assign __DOLLAR__procmux__DOLLAR__706__A[9] = __DOLLAR__procdff__DOLLAR__757__Q[9];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__A[9] = __DOLLAR__procdff__DOLLAR__757__Q[9];
  assign __DOLLAR__procmux__DOLLAR__674__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__674__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__674__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__674__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__674__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__674__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__674__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__674__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__674__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__674__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__674__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__674__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__674__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__674__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__674__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__674__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__677__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__677__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__677__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__677__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__677__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__677__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__677__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__677__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__677__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__677__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__677__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__677__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__677__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__677__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__677__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__677__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__680__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__680__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__680__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__680__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__680__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__680__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__680__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__680__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__680__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__680__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__680__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__680__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__680__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__680__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__680__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__680__B[9] = cfg_d[9];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__684_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__685_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[0] = cfg_a[0];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[1] = cfg_a[1];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[2] = cfg_a[2];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[3] = cfg_a[3];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[4] = cfg_a[4];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[5] = cfg_a[5];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[6] = cfg_a[6];
  assign __DOLLAR__procmux__DOLLAR__686_CMP0__A[7] = cfg_a[7];
  assign __DOLLAR__procmux__DOLLAR__689_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__689_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__690_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__690_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__691_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__691_CMP0__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__692_CMP0__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__692_CMP0__A[1] = data_in[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[0] = __DOLLAR__procmux__DOLLAR__693__Y[0];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[1] = __DOLLAR__procmux__DOLLAR__693__Y[1];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[10] = __DOLLAR__procmux__DOLLAR__693__Y[10];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[11] = __DOLLAR__procmux__DOLLAR__693__Y[11];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[12] = __DOLLAR__procmux__DOLLAR__693__Y[12];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[13] = __DOLLAR__procmux__DOLLAR__693__Y[13];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[14] = __DOLLAR__procmux__DOLLAR__693__Y[14];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[15] = __DOLLAR__procmux__DOLLAR__693__Y[15];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[2] = __DOLLAR__procmux__DOLLAR__693__Y[2];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[3] = __DOLLAR__procmux__DOLLAR__693__Y[3];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[4] = __DOLLAR__procmux__DOLLAR__693__Y[4];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[5] = __DOLLAR__procmux__DOLLAR__693__Y[5];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[6] = __DOLLAR__procmux__DOLLAR__693__Y[6];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[7] = __DOLLAR__procmux__DOLLAR__693__Y[7];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[8] = __DOLLAR__procmux__DOLLAR__693__Y[8];
  assign __DOLLAR__ternary__DOLLAR____DOT____DOT____FORWARD_SLASH__original_pe_verilator__FORWARD_SLASH__test_opt_reg_file__DOT__sv__COLON__119__DOLLAR__69__B[9] = __DOLLAR__procmux__DOLLAR__693__Y[9];
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__694_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__697_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__A[0] = mode[0];
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__A[1] = mode[1];
  assign __DOLLAR__procmux__DOLLAR__698_CMP0__A[2] = mode[2];
  assign __DOLLAR__procmux__DOLLAR__706__B[0] = __DOLLAR__procmux__DOLLAR__715__Y[0];
  assign __DOLLAR__procmux__DOLLAR__706__B[1] = __DOLLAR__procmux__DOLLAR__715__Y[1];
  assign __DOLLAR__procmux__DOLLAR__706__B[10] = __DOLLAR__procmux__DOLLAR__715__Y[10];
  assign __DOLLAR__procmux__DOLLAR__706__B[11] = __DOLLAR__procmux__DOLLAR__715__Y[11];
  assign __DOLLAR__procmux__DOLLAR__706__B[12] = __DOLLAR__procmux__DOLLAR__715__Y[12];
  assign __DOLLAR__procmux__DOLLAR__706__B[13] = __DOLLAR__procmux__DOLLAR__715__Y[13];
  assign __DOLLAR__procmux__DOLLAR__706__B[14] = __DOLLAR__procmux__DOLLAR__715__Y[14];
  assign __DOLLAR__procmux__DOLLAR__706__B[15] = __DOLLAR__procmux__DOLLAR__715__Y[15];
  assign __DOLLAR__procmux__DOLLAR__706__B[2] = __DOLLAR__procmux__DOLLAR__715__Y[2];
  assign __DOLLAR__procmux__DOLLAR__706__B[3] = __DOLLAR__procmux__DOLLAR__715__Y[3];
  assign __DOLLAR__procmux__DOLLAR__706__B[4] = __DOLLAR__procmux__DOLLAR__715__Y[4];
  assign __DOLLAR__procmux__DOLLAR__706__B[5] = __DOLLAR__procmux__DOLLAR__715__Y[5];
  assign __DOLLAR__procmux__DOLLAR__706__B[6] = __DOLLAR__procmux__DOLLAR__715__Y[6];
  assign __DOLLAR__procmux__DOLLAR__706__B[7] = __DOLLAR__procmux__DOLLAR__715__Y[7];
  assign __DOLLAR__procmux__DOLLAR__706__B[8] = __DOLLAR__procmux__DOLLAR__715__Y[8];
  assign __DOLLAR__procmux__DOLLAR__706__B[9] = __DOLLAR__procmux__DOLLAR__715__Y[9];
  assign __DOLLAR__procmux__DOLLAR__709__A[0] = data_in[0];
  assign __DOLLAR__procmux__DOLLAR__709__A[1] = data_in[1];
  assign __DOLLAR__procmux__DOLLAR__709__A[10] = data_in[10];
  assign __DOLLAR__procmux__DOLLAR__709__A[11] = data_in[11];
  assign __DOLLAR__procmux__DOLLAR__709__A[12] = data_in[12];
  assign __DOLLAR__procmux__DOLLAR__709__A[13] = data_in[13];
  assign __DOLLAR__procmux__DOLLAR__709__A[14] = data_in[14];
  assign __DOLLAR__procmux__DOLLAR__709__A[15] = data_in[15];
  assign __DOLLAR__procmux__DOLLAR__709__A[2] = data_in[2];
  assign __DOLLAR__procmux__DOLLAR__709__A[3] = data_in[3];
  assign __DOLLAR__procmux__DOLLAR__709__A[4] = data_in[4];
  assign __DOLLAR__procmux__DOLLAR__709__A[5] = data_in[5];
  assign __DOLLAR__procmux__DOLLAR__709__A[6] = data_in[6];
  assign __DOLLAR__procmux__DOLLAR__709__A[7] = data_in[7];
  assign __DOLLAR__procmux__DOLLAR__709__A[8] = data_in[8];
  assign __DOLLAR__procmux__DOLLAR__709__A[9] = data_in[9];
  assign __DOLLAR__procmux__DOLLAR__709__B[0] = val[0];
  assign __DOLLAR__procmux__DOLLAR__709__B[1] = val[1];
  assign __DOLLAR__procmux__DOLLAR__709__B[10] = val[10];
  assign __DOLLAR__procmux__DOLLAR__709__B[11] = val[11];
  assign __DOLLAR__procmux__DOLLAR__709__B[12] = val[12];
  assign __DOLLAR__procmux__DOLLAR__709__B[13] = val[13];
  assign __DOLLAR__procmux__DOLLAR__709__B[14] = val[14];
  assign __DOLLAR__procmux__DOLLAR__709__B[15] = val[15];
  assign __DOLLAR__procmux__DOLLAR__709__B[2] = val[2];
  assign __DOLLAR__procmux__DOLLAR__709__B[3] = val[3];
  assign __DOLLAR__procmux__DOLLAR__709__B[4] = val[4];
  assign __DOLLAR__procmux__DOLLAR__709__B[5] = val[5];
  assign __DOLLAR__procmux__DOLLAR__709__B[6] = val[6];
  assign __DOLLAR__procmux__DOLLAR__709__B[7] = val[7];
  assign __DOLLAR__procmux__DOLLAR__709__B[8] = val[8];
  assign __DOLLAR__procmux__DOLLAR__709__B[9] = val[9];
  assign __DOLLAR__procmux__DOLLAR__712__A[0] = __DOLLAR__procmux__DOLLAR__709__Y[0];
  assign __DOLLAR__procmux__DOLLAR__712__A[1] = __DOLLAR__procmux__DOLLAR__709__Y[1];
  assign __DOLLAR__procmux__DOLLAR__712__A[10] = __DOLLAR__procmux__DOLLAR__709__Y[10];
  assign __DOLLAR__procmux__DOLLAR__712__A[11] = __DOLLAR__procmux__DOLLAR__709__Y[11];
  assign __DOLLAR__procmux__DOLLAR__712__A[12] = __DOLLAR__procmux__DOLLAR__709__Y[12];
  assign __DOLLAR__procmux__DOLLAR__712__A[13] = __DOLLAR__procmux__DOLLAR__709__Y[13];
  assign __DOLLAR__procmux__DOLLAR__712__A[14] = __DOLLAR__procmux__DOLLAR__709__Y[14];
  assign __DOLLAR__procmux__DOLLAR__712__A[15] = __DOLLAR__procmux__DOLLAR__709__Y[15];
  assign __DOLLAR__procmux__DOLLAR__712__A[2] = __DOLLAR__procmux__DOLLAR__709__Y[2];
  assign __DOLLAR__procmux__DOLLAR__712__A[3] = __DOLLAR__procmux__DOLLAR__709__Y[3];
  assign __DOLLAR__procmux__DOLLAR__712__A[4] = __DOLLAR__procmux__DOLLAR__709__Y[4];
  assign __DOLLAR__procmux__DOLLAR__712__A[5] = __DOLLAR__procmux__DOLLAR__709__Y[5];
  assign __DOLLAR__procmux__DOLLAR__712__A[6] = __DOLLAR__procmux__DOLLAR__709__Y[6];
  assign __DOLLAR__procmux__DOLLAR__712__A[7] = __DOLLAR__procmux__DOLLAR__709__Y[7];
  assign __DOLLAR__procmux__DOLLAR__712__A[8] = __DOLLAR__procmux__DOLLAR__709__Y[8];
  assign __DOLLAR__procmux__DOLLAR__712__A[9] = __DOLLAR__procmux__DOLLAR__709__Y[9];
  assign __DOLLAR__procmux__DOLLAR__715__A[0] = __DOLLAR__procmux__DOLLAR__712__Y[0];
  assign __DOLLAR__procmux__DOLLAR__715__A[1] = __DOLLAR__procmux__DOLLAR__712__Y[1];
  assign __DOLLAR__procmux__DOLLAR__715__A[10] = __DOLLAR__procmux__DOLLAR__712__Y[10];
  assign __DOLLAR__procmux__DOLLAR__715__A[11] = __DOLLAR__procmux__DOLLAR__712__Y[11];
  assign __DOLLAR__procmux__DOLLAR__715__A[12] = __DOLLAR__procmux__DOLLAR__712__Y[12];
  assign __DOLLAR__procmux__DOLLAR__715__A[13] = __DOLLAR__procmux__DOLLAR__712__Y[13];
  assign __DOLLAR__procmux__DOLLAR__715__A[14] = __DOLLAR__procmux__DOLLAR__712__Y[14];
  assign __DOLLAR__procmux__DOLLAR__715__A[15] = __DOLLAR__procmux__DOLLAR__712__Y[15];
  assign __DOLLAR__procmux__DOLLAR__715__A[2] = __DOLLAR__procmux__DOLLAR__712__Y[2];
  assign __DOLLAR__procmux__DOLLAR__715__A[3] = __DOLLAR__procmux__DOLLAR__712__Y[3];
  assign __DOLLAR__procmux__DOLLAR__715__A[4] = __DOLLAR__procmux__DOLLAR__712__Y[4];
  assign __DOLLAR__procmux__DOLLAR__715__A[5] = __DOLLAR__procmux__DOLLAR__712__Y[5];
  assign __DOLLAR__procmux__DOLLAR__715__A[6] = __DOLLAR__procmux__DOLLAR__712__Y[6];
  assign __DOLLAR__procmux__DOLLAR__715__A[7] = __DOLLAR__procmux__DOLLAR__712__Y[7];
  assign __DOLLAR__procmux__DOLLAR__715__A[8] = __DOLLAR__procmux__DOLLAR__712__Y[8];
  assign __DOLLAR__procmux__DOLLAR__715__A[9] = __DOLLAR__procmux__DOLLAR__712__Y[9];
  assign __DOLLAR__procmux__DOLLAR__715__B[0] = cfg_d[0];
  assign __DOLLAR__procmux__DOLLAR__715__B[1] = cfg_d[1];
  assign __DOLLAR__procmux__DOLLAR__715__B[10] = cfg_d[10];
  assign __DOLLAR__procmux__DOLLAR__715__B[11] = cfg_d[11];
  assign __DOLLAR__procmux__DOLLAR__715__B[12] = cfg_d[12];
  assign __DOLLAR__procmux__DOLLAR__715__B[13] = cfg_d[13];
  assign __DOLLAR__procmux__DOLLAR__715__B[14] = cfg_d[14];
  assign __DOLLAR__procmux__DOLLAR__715__B[15] = cfg_d[15];
  assign __DOLLAR__procmux__DOLLAR__715__B[2] = cfg_d[2];
  assign __DOLLAR__procmux__DOLLAR__715__B[3] = cfg_d[3];
  assign __DOLLAR__procmux__DOLLAR__715__B[4] = cfg_d[4];
  assign __DOLLAR__procmux__DOLLAR__715__B[5] = cfg_d[5];
  assign __DOLLAR__procmux__DOLLAR__715__B[6] = cfg_d[6];
  assign __DOLLAR__procmux__DOLLAR__715__B[7] = cfg_d[7];
  assign __DOLLAR__procmux__DOLLAR__715__B[8] = cfg_d[8];
  assign __DOLLAR__procmux__DOLLAR__715__B[9] = cfg_d[9];

endmodule //test_opt_reg_file
